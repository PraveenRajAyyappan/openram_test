magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1335 -1309 8070 19691
<< locali >>
rect 6709 11329 6743 11345
rect 4262 11295 6709 11329
rect 6709 11279 6743 11295
rect 3374 10660 3408 10676
rect 3374 10610 3408 10626
rect 3967 10622 4001 10638
rect 3967 10572 4001 10588
rect 6709 9915 6743 9931
rect 3678 9881 6709 9915
rect 6709 9865 6743 9881
rect 3374 9170 3408 9186
rect 3374 9120 3408 9136
rect 3489 9170 3523 9186
rect 3489 9120 3523 9136
rect 6709 8501 6743 8517
rect 3678 8467 6709 8501
rect 6709 8451 6743 8467
rect 3422 8231 3456 8247
rect 3422 8181 3456 8197
rect 3522 7983 3556 7999
rect 3522 7933 3556 7949
rect 3842 7350 3876 7832
rect 4329 7831 4363 7847
rect 4329 7781 4363 7797
rect 3657 7316 3876 7350
rect 6709 7087 6743 7103
rect 4622 7053 6709 7087
rect 6709 7037 6743 7053
rect 4401 6380 4435 6396
rect 4401 6330 4435 6346
rect 3655 6191 3689 6207
rect 3655 6141 3689 6157
rect 3522 6067 3556 6083
rect 3522 6017 3556 6033
rect 3389 5943 3423 5959
rect 3389 5893 3423 5909
rect 6709 5673 6743 5689
rect 4588 5639 6709 5673
rect 6709 5623 6743 5639
rect 3389 5403 3423 5419
rect 3389 5353 3423 5369
rect 3522 5279 3556 5295
rect 3522 5229 3556 5245
rect 3655 5155 3689 5171
rect 3655 5105 3689 5121
rect 4185 4982 4219 4998
rect 4185 4932 4219 4948
rect 6709 4259 6743 4275
rect 4588 4225 6709 4259
rect 6709 4209 6743 4225
rect 4193 3536 4227 3552
rect 4193 3486 4227 3502
rect 3522 3363 3556 3379
rect 3522 3313 3556 3329
rect 3422 3115 3456 3131
rect 3422 3065 3456 3081
rect 6709 2845 6743 2861
rect 4704 2811 6709 2845
rect 6709 2795 6743 2811
rect 3639 2541 3824 2575
rect 3374 2176 3408 2192
rect 3639 2176 3673 2541
rect 3890 2327 3924 2343
rect 3890 2277 3924 2293
rect 3506 2142 3673 2176
rect 4561 2154 4595 2170
rect 3374 2126 3408 2142
rect 4561 2104 4595 2120
rect 6709 1431 6743 1447
rect 5072 1397 6709 1431
rect 6709 1381 6743 1397
rect 5785 724 5819 740
rect 3374 686 3408 702
rect 5785 674 5819 690
rect 3374 636 3408 652
rect 6709 17 6743 33
rect 6709 -33 6743 -17
<< viali >>
rect 6709 11295 6743 11329
rect 3374 10626 3408 10660
rect 3967 10588 4001 10622
rect 6709 9881 6743 9915
rect 3374 9136 3408 9170
rect 3489 9136 3523 9170
rect 6709 8467 6743 8501
rect 3422 8197 3456 8231
rect 3522 7949 3556 7983
rect 4329 7797 4363 7831
rect 6709 7053 6743 7087
rect 4401 6346 4435 6380
rect 3655 6157 3689 6191
rect 3522 6033 3556 6067
rect 3389 5909 3423 5943
rect 6709 5639 6743 5673
rect 3389 5369 3423 5403
rect 3522 5245 3556 5279
rect 3655 5121 3689 5155
rect 4185 4948 4219 4982
rect 6709 4225 6743 4259
rect 4193 3502 4227 3536
rect 3522 3329 3556 3363
rect 3422 3081 3456 3115
rect 6709 2811 6743 2845
rect 3890 2293 3924 2327
rect 3374 2142 3408 2176
rect 4561 2120 4595 2154
rect 6709 1397 6743 1431
rect 3374 652 3408 686
rect 5785 690 5819 724
rect 6709 -17 6743 17
<< metal1 >>
rect 6694 11286 6700 11338
rect 6752 11286 6758 11338
rect 2704 10617 2710 10669
rect 2762 10657 2768 10669
rect 3362 10660 3420 10666
rect 3362 10657 3374 10660
rect 2762 10629 3374 10657
rect 2762 10617 2768 10629
rect 3362 10626 3374 10629
rect 3408 10626 3420 10660
rect 3362 10620 3420 10626
rect 3952 10579 3958 10631
rect 4010 10579 4016 10631
rect 6694 9872 6700 9924
rect 6752 9872 6758 9924
rect 2620 9127 2626 9179
rect 2678 9167 2684 9179
rect 3362 9170 3420 9176
rect 3362 9167 3374 9170
rect 2678 9139 3374 9167
rect 2678 9127 2684 9139
rect 3362 9136 3374 9139
rect 3408 9136 3420 9170
rect 3362 9130 3420 9136
rect 3474 9127 3480 9179
rect 3532 9127 3538 9179
rect 6694 8458 6700 8510
rect 6752 8458 6758 8510
rect 2788 8188 2794 8240
rect 2846 8228 2852 8240
rect 3410 8231 3468 8237
rect 3410 8228 3422 8231
rect 2846 8200 3422 8228
rect 2846 8188 2852 8200
rect 3410 8197 3422 8200
rect 3456 8197 3468 8231
rect 3410 8191 3468 8197
rect 2620 7940 2626 7992
rect 2678 7980 2684 7992
rect 3510 7983 3568 7989
rect 3510 7980 3522 7983
rect 2678 7952 3522 7980
rect 2678 7940 2684 7952
rect 3510 7949 3522 7952
rect 3556 7949 3568 7983
rect 3510 7943 3568 7949
rect 4314 7788 4320 7840
rect 4372 7788 4378 7840
rect 6694 7044 6700 7096
rect 6752 7044 6758 7096
rect 4386 6337 4392 6389
rect 4444 6337 4450 6389
rect 2704 6148 2710 6200
rect 2762 6188 2768 6200
rect 3643 6191 3701 6197
rect 3643 6188 3655 6191
rect 2762 6160 3655 6188
rect 2762 6148 2768 6160
rect 3643 6157 3655 6160
rect 3689 6157 3701 6191
rect 3643 6151 3701 6157
rect 2536 6024 2542 6076
rect 2594 6064 2600 6076
rect 3510 6067 3568 6073
rect 3510 6064 3522 6067
rect 2594 6036 3522 6064
rect 2594 6024 2600 6036
rect 3510 6033 3522 6036
rect 3556 6033 3568 6067
rect 3510 6027 3568 6033
rect 2872 5900 2878 5952
rect 2930 5940 2936 5952
rect 3377 5943 3435 5949
rect 3377 5940 3389 5943
rect 2930 5912 3389 5940
rect 2930 5900 2936 5912
rect 3377 5909 3389 5912
rect 3423 5909 3435 5943
rect 3377 5903 3435 5909
rect 6694 5630 6700 5682
rect 6752 5630 6758 5682
rect 2620 5360 2626 5412
rect 2678 5400 2684 5412
rect 3377 5403 3435 5409
rect 3377 5400 3389 5403
rect 2678 5372 3389 5400
rect 2678 5360 2684 5372
rect 3377 5369 3389 5372
rect 3423 5369 3435 5403
rect 3377 5363 3435 5369
rect 2704 5236 2710 5288
rect 2762 5276 2768 5288
rect 3510 5279 3568 5285
rect 3510 5276 3522 5279
rect 2762 5248 3522 5276
rect 2762 5236 2768 5248
rect 3510 5245 3522 5248
rect 3556 5245 3568 5279
rect 3510 5239 3568 5245
rect 2956 5112 2962 5164
rect 3014 5152 3020 5164
rect 3643 5155 3701 5161
rect 3643 5152 3655 5155
rect 3014 5124 3655 5152
rect 3014 5112 3020 5124
rect 3643 5121 3655 5124
rect 3689 5121 3701 5155
rect 3643 5115 3701 5121
rect 4170 4939 4176 4991
rect 4228 4939 4234 4991
rect 1521 4296 1527 4348
rect 1579 4336 1585 4348
rect 2620 4336 2626 4348
rect 1579 4308 2626 4336
rect 1579 4296 1585 4308
rect 2620 4296 2626 4308
rect 2678 4296 2684 4348
rect 6694 4216 6700 4268
rect 6752 4216 6758 4268
rect 351 4136 357 4188
rect 409 4176 415 4188
rect 3040 4176 3046 4188
rect 409 4148 3046 4176
rect 409 4136 415 4148
rect 3040 4136 3046 4148
rect 3098 4136 3104 4188
rect 4178 3493 4184 3545
rect 4236 3493 4242 3545
rect 3124 3320 3130 3372
rect 3182 3360 3188 3372
rect 3510 3363 3568 3369
rect 3510 3360 3522 3363
rect 3182 3332 3522 3360
rect 3182 3320 3188 3332
rect 3510 3329 3522 3332
rect 3556 3329 3568 3363
rect 3510 3323 3568 3329
rect 3040 3072 3046 3124
rect 3098 3112 3104 3124
rect 3410 3115 3468 3121
rect 3410 3112 3422 3115
rect 3098 3084 3422 3112
rect 3098 3072 3104 3084
rect 3410 3081 3422 3084
rect 3456 3081 3468 3115
rect 3410 3075 3468 3081
rect 6694 2802 6700 2854
rect 6752 2802 6758 2854
rect 3875 2284 3881 2336
rect 3933 2284 3939 2336
rect 3040 2133 3046 2185
rect 3098 2173 3104 2185
rect 3362 2176 3420 2182
rect 3362 2173 3374 2176
rect 3098 2145 3374 2173
rect 3098 2133 3104 2145
rect 3362 2142 3374 2145
rect 3408 2142 3420 2176
rect 3362 2136 3420 2142
rect 4546 2111 4552 2163
rect 4604 2111 4610 2163
rect 6694 1388 6700 1440
rect 6752 1388 6758 1440
rect 3359 643 3365 695
rect 3417 643 3423 695
rect 5770 681 5776 733
rect 5828 681 5834 733
rect 6694 -26 6700 26
rect 6752 -26 6758 26
<< via1 >>
rect 6700 11329 6752 11338
rect 6700 11295 6709 11329
rect 6709 11295 6743 11329
rect 6743 11295 6752 11329
rect 6700 11286 6752 11295
rect 2710 10617 2762 10669
rect 3958 10622 4010 10631
rect 3958 10588 3967 10622
rect 3967 10588 4001 10622
rect 4001 10588 4010 10622
rect 3958 10579 4010 10588
rect 6700 9915 6752 9924
rect 6700 9881 6709 9915
rect 6709 9881 6743 9915
rect 6743 9881 6752 9915
rect 6700 9872 6752 9881
rect 2626 9127 2678 9179
rect 3480 9170 3532 9179
rect 3480 9136 3489 9170
rect 3489 9136 3523 9170
rect 3523 9136 3532 9170
rect 3480 9127 3532 9136
rect 6700 8501 6752 8510
rect 6700 8467 6709 8501
rect 6709 8467 6743 8501
rect 6743 8467 6752 8501
rect 6700 8458 6752 8467
rect 2794 8188 2846 8240
rect 2626 7940 2678 7992
rect 4320 7831 4372 7840
rect 4320 7797 4329 7831
rect 4329 7797 4363 7831
rect 4363 7797 4372 7831
rect 4320 7788 4372 7797
rect 6700 7087 6752 7096
rect 6700 7053 6709 7087
rect 6709 7053 6743 7087
rect 6743 7053 6752 7087
rect 6700 7044 6752 7053
rect 4392 6380 4444 6389
rect 4392 6346 4401 6380
rect 4401 6346 4435 6380
rect 4435 6346 4444 6380
rect 4392 6337 4444 6346
rect 2710 6148 2762 6200
rect 2542 6024 2594 6076
rect 2878 5900 2930 5952
rect 6700 5673 6752 5682
rect 6700 5639 6709 5673
rect 6709 5639 6743 5673
rect 6743 5639 6752 5673
rect 6700 5630 6752 5639
rect 2626 5360 2678 5412
rect 2710 5236 2762 5288
rect 2962 5112 3014 5164
rect 4176 4982 4228 4991
rect 4176 4948 4185 4982
rect 4185 4948 4219 4982
rect 4219 4948 4228 4982
rect 4176 4939 4228 4948
rect 1527 4296 1579 4348
rect 2626 4296 2678 4348
rect 6700 4259 6752 4268
rect 6700 4225 6709 4259
rect 6709 4225 6743 4259
rect 6743 4225 6752 4259
rect 6700 4216 6752 4225
rect 357 4136 409 4188
rect 3046 4136 3098 4188
rect 4184 3536 4236 3545
rect 4184 3502 4193 3536
rect 4193 3502 4227 3536
rect 4227 3502 4236 3536
rect 4184 3493 4236 3502
rect 3130 3320 3182 3372
rect 3046 3072 3098 3124
rect 6700 2845 6752 2854
rect 6700 2811 6709 2845
rect 6709 2811 6743 2845
rect 6743 2811 6752 2845
rect 6700 2802 6752 2811
rect 3881 2327 3933 2336
rect 3881 2293 3890 2327
rect 3890 2293 3924 2327
rect 3924 2293 3933 2327
rect 3881 2284 3933 2293
rect 3046 2133 3098 2185
rect 4552 2154 4604 2163
rect 4552 2120 4561 2154
rect 4561 2120 4595 2154
rect 4595 2120 4604 2154
rect 4552 2111 4604 2120
rect 6700 1431 6752 1440
rect 6700 1397 6709 1431
rect 6709 1397 6743 1431
rect 6743 1397 6752 1431
rect 6700 1388 6752 1397
rect 3365 686 3417 695
rect 3365 652 3374 686
rect 3374 652 3408 686
rect 3408 652 3417 686
rect 3365 643 3417 652
rect 5776 724 5828 733
rect 5776 690 5785 724
rect 5785 690 5819 724
rect 5819 690 5828 724
rect 5776 681 5828 690
rect 6700 17 6752 26
rect 6700 -17 6709 17
rect 6709 -17 6743 17
rect 6743 -17 6752 17
rect 6700 -26 6752 -17
<< metal2 >>
rect -57 17699 -29 17727
rect 2554 8624 2582 11352
rect 2638 9185 2666 11352
rect 2722 10675 2750 11352
rect 2710 10669 2762 10675
rect 2710 10611 2762 10617
rect 2626 9179 2678 9185
rect 2626 9121 2678 9127
rect 2540 8615 2596 8624
rect 2540 8550 2596 8559
rect 1539 4354 1567 6401
rect 2554 6082 2582 8550
rect 2638 7998 2666 9121
rect 2626 7992 2678 7998
rect 2626 7934 2678 7940
rect 2542 6076 2594 6082
rect 2542 6018 2594 6024
rect 1527 4348 1579 4354
rect 1527 4290 1579 4296
rect 357 4188 409 4194
rect 357 4130 409 4136
rect 369 2828 397 4130
rect 2350 2353 2406 2362
rect 137 2238 203 2290
rect 2350 2288 2406 2297
rect 1844 1971 1900 1980
rect 1844 1906 1900 1915
rect 1844 913 1900 922
rect 1844 848 1900 857
rect 137 538 203 590
rect 2554 0 2582 6018
rect 2638 5418 2666 7934
rect 2722 6206 2750 10611
rect 2806 8246 2834 11352
rect 2794 8240 2846 8246
rect 2794 8182 2846 8188
rect 2710 6200 2762 6206
rect 2710 6142 2762 6148
rect 2626 5412 2678 5418
rect 2626 5354 2678 5360
rect 2638 4354 2666 5354
rect 2722 5294 2750 6142
rect 2710 5288 2762 5294
rect 2710 5230 2762 5236
rect 2626 4348 2678 4354
rect 2626 4290 2678 4296
rect 2638 0 2666 4290
rect 2722 1608 2750 5230
rect 2806 3556 2834 8182
rect 2890 5958 2918 11352
rect 2878 5952 2930 5958
rect 2878 5894 2930 5900
rect 2792 3547 2848 3556
rect 2792 3482 2848 3491
rect 2708 1599 2764 1608
rect 2708 1534 2764 1543
rect 2722 0 2750 1534
rect 2806 0 2834 3482
rect 2890 1980 2918 5894
rect 2974 5170 3002 11352
rect 2962 5164 3014 5170
rect 2962 5106 3014 5112
rect 2974 2362 3002 5106
rect 3058 4194 3086 11352
rect 3046 4188 3098 4194
rect 3046 4130 3098 4136
rect 3058 3130 3086 4130
rect 3142 3378 3170 11352
rect 6698 11340 6754 11349
rect 6698 11275 6754 11284
rect 3958 10631 4010 10637
rect 4010 10591 6810 10619
rect 3958 10573 4010 10579
rect 6698 9926 6754 9935
rect 6698 9861 6754 9870
rect 3480 9179 3532 9185
rect 3480 9121 3532 9127
rect 3492 8624 3520 9121
rect 3478 8615 3534 8624
rect 3478 8550 3534 8559
rect 6698 8512 6754 8521
rect 6698 8447 6754 8456
rect 4320 7840 4372 7846
rect 4372 7800 6810 7828
rect 4320 7782 4372 7788
rect 6698 7098 6754 7107
rect 6698 7033 6754 7042
rect 4392 6389 4444 6395
rect 4444 6349 6810 6377
rect 4392 6331 4444 6337
rect 6698 5684 6754 5693
rect 6698 5619 6754 5628
rect 4176 4991 4228 4997
rect 4228 4951 6810 4979
rect 4176 4933 4228 4939
rect 6698 4270 6754 4279
rect 6698 4205 6754 4214
rect 4182 3547 4238 3556
rect 4182 3482 4238 3491
rect 3130 3372 3182 3378
rect 3130 3314 3182 3320
rect 3046 3124 3098 3130
rect 3046 3066 3098 3072
rect 2960 2353 3016 2362
rect 2960 2288 3016 2297
rect 2876 1971 2932 1980
rect 2876 1906 2932 1915
rect 2890 0 2918 1906
rect 2974 0 3002 2288
rect 3058 2191 3086 3066
rect 3142 2347 3170 3314
rect 6698 2856 6754 2865
rect 6698 2791 6754 2800
rect 3128 2338 3184 2347
rect 3128 2273 3184 2282
rect 3879 2338 3935 2347
rect 3879 2273 3935 2282
rect 3046 2185 3098 2191
rect 3046 2127 3098 2133
rect 3058 178 3086 2127
rect 3142 922 3170 2273
rect 4552 2163 4604 2169
rect 4552 2105 4604 2111
rect 4564 1608 4592 2105
rect 4550 1599 4606 1608
rect 4550 1534 4606 1543
rect 6698 1442 6754 1451
rect 6698 1377 6754 1386
rect 3128 913 3184 922
rect 3128 848 3184 857
rect 3044 169 3100 178
rect 3044 104 3100 113
rect 3058 0 3086 104
rect 3142 0 3170 848
rect 5776 733 5828 739
rect 3365 695 3417 701
rect 5828 693 6810 721
rect 5776 675 5828 681
rect 3365 637 3417 643
rect 5788 178 5816 675
rect 5774 169 5830 178
rect 5774 104 5830 113
rect 6698 28 6754 37
rect 6698 -37 6754 -28
<< via2 >>
rect 2540 8559 2596 8615
rect 2350 2297 2406 2353
rect 1844 1915 1900 1971
rect 1844 857 1900 913
rect 2792 3491 2848 3547
rect 2708 1543 2764 1599
rect 6698 11338 6754 11340
rect 6698 11286 6700 11338
rect 6700 11286 6752 11338
rect 6752 11286 6754 11338
rect 6698 11284 6754 11286
rect 6698 9924 6754 9926
rect 6698 9872 6700 9924
rect 6700 9872 6752 9924
rect 6752 9872 6754 9924
rect 6698 9870 6754 9872
rect 3478 8559 3534 8615
rect 6698 8510 6754 8512
rect 6698 8458 6700 8510
rect 6700 8458 6752 8510
rect 6752 8458 6754 8510
rect 6698 8456 6754 8458
rect 6698 7096 6754 7098
rect 6698 7044 6700 7096
rect 6700 7044 6752 7096
rect 6752 7044 6754 7096
rect 6698 7042 6754 7044
rect 6698 5682 6754 5684
rect 6698 5630 6700 5682
rect 6700 5630 6752 5682
rect 6752 5630 6754 5682
rect 6698 5628 6754 5630
rect 6698 4268 6754 4270
rect 6698 4216 6700 4268
rect 6700 4216 6752 4268
rect 6752 4216 6754 4268
rect 6698 4214 6754 4216
rect 4182 3545 4238 3547
rect 4182 3493 4184 3545
rect 4184 3493 4236 3545
rect 4236 3493 4238 3545
rect 4182 3491 4238 3493
rect 2960 2297 3016 2353
rect 2876 1915 2932 1971
rect 6698 2854 6754 2856
rect 6698 2802 6700 2854
rect 6700 2802 6752 2854
rect 6752 2802 6754 2854
rect 6698 2800 6754 2802
rect 3128 2282 3184 2338
rect 3879 2336 3935 2338
rect 3879 2284 3881 2336
rect 3881 2284 3933 2336
rect 3933 2284 3935 2336
rect 3879 2282 3935 2284
rect 4550 1543 4606 1599
rect 6698 1440 6754 1442
rect 6698 1388 6700 1440
rect 6700 1388 6752 1440
rect 6752 1388 6754 1440
rect 6698 1386 6754 1388
rect 3128 857 3184 913
rect 3044 113 3100 169
rect 5774 113 5830 169
rect 6698 26 6754 28
rect 6698 -26 6700 26
rect 6700 -26 6752 26
rect 6752 -26 6754 26
rect 6698 -28 6754 -26
<< metal3 >>
rect 607 18333 705 18431
rect 1343 18333 1441 18431
rect 607 16919 705 17017
rect 1343 16919 1441 17017
rect 607 15505 705 15603
rect 1343 15505 1441 15603
rect 607 14091 705 14189
rect 1343 14091 1441 14189
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 6677 11340 6775 11361
rect 6677 11284 6698 11340
rect 6754 11284 6775 11340
rect 6677 11263 6775 11284
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 6677 9926 6775 9947
rect 6677 9870 6698 9926
rect 6754 9870 6775 9926
rect 6677 9849 6775 9870
rect 2535 8617 2601 8620
rect 3473 8617 3539 8620
rect 2535 8615 3539 8617
rect 2535 8559 2540 8615
rect 2596 8559 3478 8615
rect 3534 8559 3539 8615
rect 2535 8557 3539 8559
rect 2535 8554 2601 8557
rect 3473 8554 3539 8557
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 6677 8512 6775 8533
rect 6677 8456 6698 8512
rect 6754 8456 6775 8512
rect 6677 8435 6775 8456
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 6677 7098 6775 7119
rect 6677 7042 6698 7098
rect 6754 7042 6775 7098
rect 6677 7021 6775 7042
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 6677 5684 6775 5705
rect 6677 5628 6698 5684
rect 6754 5628 6775 5684
rect 6677 5607 6775 5628
rect 6677 4270 6775 4291
rect 6677 4214 6698 4270
rect 6754 4214 6775 4270
rect 6677 4193 6775 4214
rect 2787 3549 2853 3552
rect 4177 3549 4243 3552
rect 2787 3547 4243 3549
rect 2787 3491 2792 3547
rect 2848 3491 4182 3547
rect 4238 3491 4243 3547
rect 2787 3489 4243 3491
rect 2787 3486 2853 3489
rect 4177 3486 4243 3489
rect -49 2779 49 2877
rect 6677 2856 6775 2877
rect 6677 2800 6698 2856
rect 6754 2800 6775 2856
rect 6677 2779 6775 2800
rect 2345 2355 2411 2358
rect 2955 2355 3021 2358
rect 2345 2353 3021 2355
rect 2345 2297 2350 2353
rect 2406 2297 2960 2353
rect 3016 2297 3021 2353
rect 2345 2295 3021 2297
rect 2345 2292 2411 2295
rect 2955 2292 3021 2295
rect 3123 2340 3189 2343
rect 3874 2340 3940 2343
rect 3123 2338 3940 2340
rect 3123 2282 3128 2338
rect 3184 2282 3879 2338
rect 3935 2282 3940 2338
rect 3123 2280 3940 2282
rect 3123 2277 3189 2280
rect 3874 2277 3940 2280
rect 1839 1973 1905 1976
rect 2871 1973 2937 1976
rect 1839 1971 2937 1973
rect 1839 1915 1844 1971
rect 1900 1915 2876 1971
rect 2932 1915 2937 1971
rect 1839 1913 2937 1915
rect 1839 1910 1905 1913
rect 2871 1910 2937 1913
rect 2703 1601 2769 1604
rect 4545 1601 4611 1604
rect 2703 1599 4611 1601
rect 2703 1543 2708 1599
rect 2764 1543 4550 1599
rect 4606 1543 4611 1599
rect 2703 1541 4611 1543
rect 2703 1538 2769 1541
rect 4545 1538 4611 1541
rect -49 1365 49 1463
rect 6677 1442 6775 1463
rect 6677 1386 6698 1442
rect 6754 1386 6775 1442
rect 6677 1365 6775 1386
rect 1839 915 1905 918
rect 3123 915 3189 918
rect 1839 913 3189 915
rect 1839 857 1844 913
rect 1900 857 3128 913
rect 3184 857 3189 913
rect 1839 855 3189 857
rect 1839 852 1905 855
rect 3123 852 3189 855
rect 3039 171 3105 174
rect 5769 171 5835 174
rect 3039 169 5835 171
rect 3039 113 3044 169
rect 3100 113 5774 169
rect 5830 113 5835 169
rect 3039 111 5835 113
rect 3039 108 3105 111
rect 5769 108 5835 111
rect -49 -49 49 49
rect 6677 28 6775 49
rect 6677 -28 6698 28
rect 6754 -28 6775 28
rect 6677 -49 6775 -28
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 6693 0 1 11275
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 6694 0 1 11280
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 6697 0 1 11279
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 6693 0 1 9861
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 6694 0 1 9866
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 6697 0 1 9865
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 6693 0 1 8447
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 6694 0 1 8452
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 6697 0 1 8451
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 6693 0 1 9861
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 6694 0 1 9866
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 6697 0 1 9865
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 6693 0 1 8447
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 6694 0 1 8452
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 6697 0 1 8451
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 6693 0 1 7033
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 6694 0 1 7038
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 6697 0 1 7037
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 6693 0 1 5619
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 6694 0 1 5624
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 6697 0 1 5623
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 6693 0 1 7033
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 6694 0 1 7038
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 6697 0 1 7037
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 6693 0 1 5619
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 6694 0 1 5624
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 6697 0 1 5623
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 6693 0 1 4205
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 6694 0 1 4210
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 6697 0 1 4209
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 6693 0 1 2791
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 6694 0 1 2796
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 6697 0 1 2795
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 6693 0 1 4205
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 6694 0 1 4210
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 6697 0 1 4209
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 6693 0 1 2791
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 6694 0 1 2796
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1634918361
transform 1 0 6697 0 1 2795
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 6693 0 1 1377
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 6694 0 1 1382
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1634918361
transform 1 0 6697 0 1 1381
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 6693 0 1 -37
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 6694 0 1 -32
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1634918361
transform 1 0 6697 0 1 -33
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 6693 0 1 1377
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 6694 0 1 1382
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1634918361
transform 1 0 6697 0 1 1381
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1634918361
transform 1 0 4178 0 1 3487
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1634918361
transform 1 0 4181 0 1 3486
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 4177 0 1 3482
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1634918361
transform 1 0 4178 0 1 3487
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1634918361
transform 1 0 4181 0 1 3486
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1634918361
transform 1 0 2787 0 1 3482
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1634918361
transform 1 0 3510 0 1 3313
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1634918361
transform 1 0 3124 0 1 3314
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1634918361
transform 1 0 3410 0 1 3065
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1634918361
transform 1 0 3040 0 1 3066
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1634918361
transform 1 0 4546 0 1 2105
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1634918361
transform 1 0 4549 0 1 2104
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1634918361
transform 1 0 2703 0 1 1534
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1634918361
transform 1 0 4545 0 1 1534
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1634918361
transform 1 0 3874 0 1 2273
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1634918361
transform 1 0 3875 0 1 2278
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1634918361
transform 1 0 3878 0 1 2277
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1634918361
transform 1 0 3874 0 1 2273
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1634918361
transform 1 0 3875 0 1 2278
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1634918361
transform 1 0 3878 0 1 2277
box 0 0 1 1
use contact_29  contact_29_3
timestamp 1634918361
transform 1 0 3123 0 1 2273
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1634918361
transform 1 0 3362 0 1 2126
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1634918361
transform 1 0 3040 0 1 2127
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1634918361
transform 1 0 5770 0 1 675
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1634918361
transform 1 0 5773 0 1 674
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1634918361
transform 1 0 5770 0 1 675
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1634918361
transform 1 0 5773 0 1 674
box 0 0 1 1
use contact_29  contact_29_4
timestamp 1634918361
transform 1 0 3039 0 1 104
box 0 0 1 1
use contact_29  contact_29_5
timestamp 1634918361
transform 1 0 5769 0 1 104
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1634918361
transform 1 0 3359 0 1 637
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1634918361
transform 1 0 3362 0 1 636
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1634918361
transform 1 0 4314 0 1 7782
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1634918361
transform 1 0 4317 0 1 7781
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1634918361
transform 1 0 3510 0 1 7933
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1634918361
transform 1 0 2620 0 1 7934
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1634918361
transform 1 0 3410 0 1 8181
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1634918361
transform 1 0 2788 0 1 8182
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1634918361
transform 1 0 2620 0 1 4290
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1634918361
transform 1 0 1521 0 1 4290
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1634918361
transform 1 0 4170 0 1 4933
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1634918361
transform 1 0 4173 0 1 4932
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1634918361
transform 1 0 3643 0 1 5105
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1634918361
transform 1 0 2956 0 1 5106
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1634918361
transform 1 0 3510 0 1 5229
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1634918361
transform 1 0 2704 0 1 5230
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1634918361
transform 1 0 3377 0 1 5353
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1634918361
transform 1 0 2620 0 1 5354
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1634918361
transform 1 0 4386 0 1 6331
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1634918361
transform 1 0 4389 0 1 6330
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1634918361
transform 1 0 3643 0 1 6141
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1634918361
transform 1 0 2704 0 1 6142
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1634918361
transform 1 0 3510 0 1 6017
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1634918361
transform 1 0 2536 0 1 6018
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1634918361
transform 1 0 3377 0 1 5893
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1634918361
transform 1 0 2872 0 1 5894
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1634918361
transform 1 0 3362 0 1 9120
box 0 0 1 1
use contact_19  contact_19_40
timestamp 1634918361
transform 1 0 2620 0 1 9121
box 0 0 1 1
use contact_19  contact_19_41
timestamp 1634918361
transform 1 0 3474 0 1 9121
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1634918361
transform 1 0 3477 0 1 9120
box 0 0 1 1
use contact_29  contact_29_6
timestamp 1634918361
transform 1 0 2535 0 1 8550
box 0 0 1 1
use contact_29  contact_29_7
timestamp 1634918361
transform 1 0 3473 0 1 8550
box 0 0 1 1
use contact_19  contact_19_42
timestamp 1634918361
transform 1 0 3952 0 1 10573
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1634918361
transform 1 0 3955 0 1 10572
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1634918361
transform 1 0 3362 0 1 10610
box 0 0 1 1
use contact_19  contact_19_43
timestamp 1634918361
transform 1 0 2704 0 1 10611
box 0 0 1 1
use contact_19  contact_19_44
timestamp 1634918361
transform 1 0 3040 0 1 4130
box 0 0 1 1
use contact_19  contact_19_45
timestamp 1634918361
transform 1 0 351 0 1 4130
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1634918361
transform 1 0 2345 0 1 2288
box 0 0 1 1
use contact_29  contact_29_8
timestamp 1634918361
transform 1 0 2955 0 1 2288
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1634918361
transform 1 0 1839 0 1 1906
box 0 0 1 1
use contact_29  contact_29_9
timestamp 1634918361
transform 1 0 2871 0 1 1906
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1634918361
transform 1 0 1839 0 1 848
box 0 0 1 1
use contact_29  contact_29_10
timestamp 1634918361
transform 1 0 3123 0 1 848
box 0 0 1 1
use pdriver_5  pdriver_5_0
timestamp 1634918361
transform 1 0 3778 0 -1 8484
box -36 -17 880 1471
use pnand2_1  pnand2_1_0
timestamp 1634918361
transform 1 0 3310 0 -1 8484
box -36 -17 504 1471
use delay_chain  delay_chain_0
timestamp 1634918361
transform 1 0 0 0 -1 18382
box -75 -49 1876 12783
use pand3_0  pand3_0_0
timestamp 1634918361
transform 1 0 3310 0 -1 5656
box -36 -17 1314 1471
use pand3  pand3_0
timestamp 1634918361
transform 1 0 3310 0 1 5656
box -36 -17 1746 1471
use pinv_10  pinv_10_0
timestamp 1634918361
transform 1 0 3310 0 1 8484
box -36 -17 404 1471
use pdriver_2  pdriver_2_0
timestamp 1634918361
transform 1 0 3310 0 -1 11312
box -36 -17 988 1471
use pand2_0  pand2_0_0
timestamp 1634918361
transform 1 0 3310 0 1 2828
box -36 -17 1430 1471
use pand2_0  pand2_0_1
timestamp 1634918361
transform 1 0 3678 0 -1 2828
box -36 -17 1430 1471
use pinv_10  pinv_10_1
timestamp 1634918361
transform 1 0 3310 0 -1 2828
box -36 -17 404 1471
use pdriver_1  pdriver_1_0
timestamp 1634918361
transform 1 0 3310 0 1 0
box -36 -17 3452 1471
use dff_buf_array  dff_buf_array_0
timestamp 1634918361
transform 1 0 0 0 1 0
box -49 -49 2590 2877
<< labels >>
rlabel metal2 s 137 538 203 590 4 csb
port 1 nsew
rlabel metal2 s 137 2238 203 2290 4 web
port 2 nsew
rlabel metal2 s 3984 10591 6810 10619 4 wl_en
port 3 nsew
rlabel metal2 s 4418 6349 6810 6377 4 w_en
port 4 nsew
rlabel metal2 s 4202 4951 6810 4979 4 s_en
port 5 nsew
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
port 6 nsew
rlabel metal2 s 4346 7800 6810 7828 4 p_en_bar
port 7 nsew
rlabel metal2 s 3377 655 3405 683 4 clk
port 8 nsew
rlabel metal2 s 5802 693 6810 721 4 clk_buf
port 9 nsew
rlabel metal3 s 1343 5607 1441 5705 4 vdd
port 10 nsew
rlabel metal3 s 1343 11263 1441 11361 4 vdd
port 10 nsew
rlabel metal3 s 1343 14091 1441 14189 4 vdd
port 10 nsew
rlabel metal3 s 607 14091 705 14189 4 vdd
port 10 nsew
rlabel metal3 s 607 11263 705 11361 4 vdd
port 10 nsew
rlabel metal3 s 6677 7021 6775 7119 4 vdd
port 10 nsew
rlabel metal3 s 6677 9849 6775 9947 4 vdd
port 10 nsew
rlabel metal3 s 1343 16919 1441 17017 4 vdd
port 10 nsew
rlabel metal3 s 607 8435 705 8533 4 vdd
port 10 nsew
rlabel metal3 s 607 5607 705 5705 4 vdd
port 10 nsew
rlabel metal3 s 6677 1365 6775 1463 4 vdd
port 10 nsew
rlabel metal3 s 607 16919 705 17017 4 vdd
port 10 nsew
rlabel metal3 s 6677 4193 6775 4291 4 vdd
port 10 nsew
rlabel metal3 s -49 1365 49 1463 4 vdd
port 10 nsew
rlabel metal3 s 1343 8435 1441 8533 4 vdd
port 10 nsew
rlabel metal3 s 607 15505 705 15603 4 gnd
port 11 nsew
rlabel metal3 s 1343 15505 1441 15603 4 gnd
port 11 nsew
rlabel metal3 s 6677 -49 6775 49 4 gnd
port 11 nsew
rlabel metal3 s 6677 8435 6775 8533 4 gnd
port 11 nsew
rlabel metal3 s 607 18333 705 18431 4 gnd
port 11 nsew
rlabel metal3 s 607 7021 705 7119 4 gnd
port 11 nsew
rlabel metal3 s 1343 18333 1441 18431 4 gnd
port 11 nsew
rlabel metal3 s 1343 9849 1441 9947 4 gnd
port 11 nsew
rlabel metal3 s 6677 11263 6775 11361 4 gnd
port 11 nsew
rlabel metal3 s 607 9849 705 9947 4 gnd
port 11 nsew
rlabel metal3 s 6677 2779 6775 2877 4 gnd
port 11 nsew
rlabel metal3 s -49 2779 49 2877 4 gnd
port 11 nsew
rlabel metal3 s 6677 5607 6775 5705 4 gnd
port 11 nsew
rlabel metal3 s 607 12677 705 12775 4 gnd
port 11 nsew
rlabel metal3 s -49 -49 49 49 4 gnd
port 11 nsew
rlabel metal3 s 1343 7021 1441 7119 4 gnd
port 11 nsew
rlabel metal3 s 1343 12677 1441 12775 4 gnd
port 11 nsew
<< properties >>
string FIXED_BBOX 6693 -37 6759 0
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1053496
string GDS_START 1032652
<< end >>
