magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1302 -1365 6294 7685
<< metal1 >>
rect 78 0 114 6320
rect 150 0 186 6320
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 79 258 711
rect 294 0 330 6320
rect 366 0 402 6320
rect 846 0 882 6320
rect 918 0 954 6320
rect 990 5609 1026 6241
rect 990 4819 1026 5451
rect 990 4029 1026 4661
rect 990 3239 1026 3871
rect 990 2449 1026 3081
rect 990 1659 1026 2291
rect 990 869 1026 1501
rect 990 79 1026 711
rect 1062 0 1098 6320
rect 1134 0 1170 6320
rect 1326 0 1362 6320
rect 1398 0 1434 6320
rect 1470 5609 1506 6241
rect 1470 4819 1506 5451
rect 1470 4029 1506 4661
rect 1470 3239 1506 3871
rect 1470 2449 1506 3081
rect 1470 1659 1506 2291
rect 1470 869 1506 1501
rect 1470 79 1506 711
rect 1542 0 1578 6320
rect 1614 0 1650 6320
rect 2094 0 2130 6320
rect 2166 0 2202 6320
rect 2238 5609 2274 6241
rect 2238 4819 2274 5451
rect 2238 4029 2274 4661
rect 2238 3239 2274 3871
rect 2238 2449 2274 3081
rect 2238 1659 2274 2291
rect 2238 869 2274 1501
rect 2238 79 2274 711
rect 2310 0 2346 6320
rect 2382 0 2418 6320
rect 2574 0 2610 6320
rect 2646 0 2682 6320
rect 2718 5609 2754 6241
rect 2718 4819 2754 5451
rect 2718 4029 2754 4661
rect 2718 3239 2754 3871
rect 2718 2449 2754 3081
rect 2718 1659 2754 2291
rect 2718 869 2754 1501
rect 2718 79 2754 711
rect 2790 0 2826 6320
rect 2862 0 2898 6320
rect 3342 0 3378 6320
rect 3414 0 3450 6320
rect 3486 5609 3522 6241
rect 3486 4819 3522 5451
rect 3486 4029 3522 4661
rect 3486 3239 3522 3871
rect 3486 2449 3522 3081
rect 3486 1659 3522 2291
rect 3486 869 3522 1501
rect 3486 79 3522 711
rect 3558 0 3594 6320
rect 3630 0 3666 6320
rect 3822 0 3858 6320
rect 3894 0 3930 6320
rect 3966 5609 4002 6241
rect 3966 4819 4002 5451
rect 3966 4029 4002 4661
rect 3966 3239 4002 3871
rect 3966 2449 4002 3081
rect 3966 1659 4002 2291
rect 3966 869 4002 1501
rect 3966 79 4002 711
rect 4038 0 4074 6320
rect 4110 0 4146 6320
rect 4590 0 4626 6320
rect 4662 0 4698 6320
rect 4734 5609 4770 6241
rect 4734 4819 4770 5451
rect 4734 4029 4770 4661
rect 4734 3239 4770 3871
rect 4734 2449 4770 3081
rect 4734 1659 4770 2291
rect 4734 869 4770 1501
rect 4734 79 4770 711
rect 4806 0 4842 6320
rect 4878 0 4914 6320
<< metal2 >>
rect 186 6265 294 6375
rect 954 6265 1062 6375
rect 1434 6265 1542 6375
rect 2202 6265 2310 6375
rect 2682 6265 2790 6375
rect 3450 6265 3558 6375
rect 3930 6265 4038 6375
rect 4698 6265 4806 6375
rect 0 6169 4992 6217
rect 186 6045 294 6121
rect 954 6045 1062 6121
rect 1434 6045 1542 6121
rect 2202 6045 2310 6121
rect 2682 6045 2790 6121
rect 3450 6045 3558 6121
rect 3930 6045 4038 6121
rect 4698 6045 4806 6121
rect 0 5949 4992 5997
rect 0 5853 4992 5901
rect 186 5729 294 5805
rect 954 5729 1062 5805
rect 1434 5729 1542 5805
rect 2202 5729 2310 5805
rect 2682 5729 2790 5805
rect 3450 5729 3558 5805
rect 3930 5729 4038 5805
rect 4698 5729 4806 5805
rect 0 5633 4992 5681
rect 186 5475 294 5585
rect 954 5475 1062 5585
rect 1434 5475 1542 5585
rect 2202 5475 2310 5585
rect 2682 5475 2790 5585
rect 3450 5475 3558 5585
rect 3930 5475 4038 5585
rect 4698 5475 4806 5585
rect 0 5379 4992 5427
rect 186 5255 294 5331
rect 954 5255 1062 5331
rect 1434 5255 1542 5331
rect 2202 5255 2310 5331
rect 2682 5255 2790 5331
rect 3450 5255 3558 5331
rect 3930 5255 4038 5331
rect 4698 5255 4806 5331
rect 0 5159 4992 5207
rect 0 5063 4992 5111
rect 186 4939 294 5015
rect 954 4939 1062 5015
rect 1434 4939 1542 5015
rect 2202 4939 2310 5015
rect 2682 4939 2790 5015
rect 3450 4939 3558 5015
rect 3930 4939 4038 5015
rect 4698 4939 4806 5015
rect 0 4843 4992 4891
rect 186 4685 294 4795
rect 954 4685 1062 4795
rect 1434 4685 1542 4795
rect 2202 4685 2310 4795
rect 2682 4685 2790 4795
rect 3450 4685 3558 4795
rect 3930 4685 4038 4795
rect 4698 4685 4806 4795
rect 0 4589 4992 4637
rect 186 4465 294 4541
rect 954 4465 1062 4541
rect 1434 4465 1542 4541
rect 2202 4465 2310 4541
rect 2682 4465 2790 4541
rect 3450 4465 3558 4541
rect 3930 4465 4038 4541
rect 4698 4465 4806 4541
rect 0 4369 4992 4417
rect 0 4273 4992 4321
rect 186 4149 294 4225
rect 954 4149 1062 4225
rect 1434 4149 1542 4225
rect 2202 4149 2310 4225
rect 2682 4149 2790 4225
rect 3450 4149 3558 4225
rect 3930 4149 4038 4225
rect 4698 4149 4806 4225
rect 0 4053 4992 4101
rect 186 3895 294 4005
rect 954 3895 1062 4005
rect 1434 3895 1542 4005
rect 2202 3895 2310 4005
rect 2682 3895 2790 4005
rect 3450 3895 3558 4005
rect 3930 3895 4038 4005
rect 4698 3895 4806 4005
rect 0 3799 4992 3847
rect 186 3675 294 3751
rect 954 3675 1062 3751
rect 1434 3675 1542 3751
rect 2202 3675 2310 3751
rect 2682 3675 2790 3751
rect 3450 3675 3558 3751
rect 3930 3675 4038 3751
rect 4698 3675 4806 3751
rect 0 3579 4992 3627
rect 0 3483 4992 3531
rect 186 3359 294 3435
rect 954 3359 1062 3435
rect 1434 3359 1542 3435
rect 2202 3359 2310 3435
rect 2682 3359 2790 3435
rect 3450 3359 3558 3435
rect 3930 3359 4038 3435
rect 4698 3359 4806 3435
rect 0 3263 4992 3311
rect 186 3105 294 3215
rect 954 3105 1062 3215
rect 1434 3105 1542 3215
rect 2202 3105 2310 3215
rect 2682 3105 2790 3215
rect 3450 3105 3558 3215
rect 3930 3105 4038 3215
rect 4698 3105 4806 3215
rect 0 3009 4992 3057
rect 186 2885 294 2961
rect 954 2885 1062 2961
rect 1434 2885 1542 2961
rect 2202 2885 2310 2961
rect 2682 2885 2790 2961
rect 3450 2885 3558 2961
rect 3930 2885 4038 2961
rect 4698 2885 4806 2961
rect 0 2789 4992 2837
rect 0 2693 4992 2741
rect 186 2569 294 2645
rect 954 2569 1062 2645
rect 1434 2569 1542 2645
rect 2202 2569 2310 2645
rect 2682 2569 2790 2645
rect 3450 2569 3558 2645
rect 3930 2569 4038 2645
rect 4698 2569 4806 2645
rect 0 2473 4992 2521
rect 186 2315 294 2425
rect 954 2315 1062 2425
rect 1434 2315 1542 2425
rect 2202 2315 2310 2425
rect 2682 2315 2790 2425
rect 3450 2315 3558 2425
rect 3930 2315 4038 2425
rect 4698 2315 4806 2425
rect 0 2219 4992 2267
rect 186 2095 294 2171
rect 954 2095 1062 2171
rect 1434 2095 1542 2171
rect 2202 2095 2310 2171
rect 2682 2095 2790 2171
rect 3450 2095 3558 2171
rect 3930 2095 4038 2171
rect 4698 2095 4806 2171
rect 0 1999 4992 2047
rect 0 1903 4992 1951
rect 186 1779 294 1855
rect 954 1779 1062 1855
rect 1434 1779 1542 1855
rect 2202 1779 2310 1855
rect 2682 1779 2790 1855
rect 3450 1779 3558 1855
rect 3930 1779 4038 1855
rect 4698 1779 4806 1855
rect 0 1683 4992 1731
rect 186 1525 294 1635
rect 954 1525 1062 1635
rect 1434 1525 1542 1635
rect 2202 1525 2310 1635
rect 2682 1525 2790 1635
rect 3450 1525 3558 1635
rect 3930 1525 4038 1635
rect 4698 1525 4806 1635
rect 0 1429 4992 1477
rect 186 1305 294 1381
rect 954 1305 1062 1381
rect 1434 1305 1542 1381
rect 2202 1305 2310 1381
rect 2682 1305 2790 1381
rect 3450 1305 3558 1381
rect 3930 1305 4038 1381
rect 4698 1305 4806 1381
rect 0 1209 4992 1257
rect 0 1113 4992 1161
rect 186 989 294 1065
rect 954 989 1062 1065
rect 1434 989 1542 1065
rect 2202 989 2310 1065
rect 2682 989 2790 1065
rect 3450 989 3558 1065
rect 3930 989 4038 1065
rect 4698 989 4806 1065
rect 0 893 4992 941
rect 186 735 294 845
rect 954 735 1062 845
rect 1434 735 1542 845
rect 2202 735 2310 845
rect 2682 735 2790 845
rect 3450 735 3558 845
rect 3930 735 4038 845
rect 4698 735 4806 845
rect 0 639 4992 687
rect 186 515 294 591
rect 954 515 1062 591
rect 1434 515 1542 591
rect 2202 515 2310 591
rect 2682 515 2790 591
rect 3450 515 3558 591
rect 3930 515 4038 591
rect 4698 515 4806 591
rect 0 419 4992 467
rect 0 323 4992 371
rect 186 199 294 275
rect 954 199 1062 275
rect 1434 199 1542 275
rect 2202 199 2310 275
rect 2682 199 2790 275
rect 3450 199 3558 275
rect 3930 199 4038 275
rect 4698 199 4806 275
rect 0 103 4992 151
rect 186 -55 294 55
rect 954 -55 1062 55
rect 1434 -55 1542 55
rect 2202 -55 2310 55
rect 2682 -55 2790 55
rect 3450 -55 3558 55
rect 3930 -55 4038 55
rect 4698 -55 4806 55
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_0
timestamp 1634918361
transform -1 0 4992 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1
timestamp 1634918361
transform -1 0 4992 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2
timestamp 1634918361
transform -1 0 4992 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_3
timestamp 1634918361
transform -1 0 4992 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_4
timestamp 1634918361
transform -1 0 4992 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_5
timestamp 1634918361
transform -1 0 4992 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_6
timestamp 1634918361
transform -1 0 4992 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_7
timestamp 1634918361
transform -1 0 4992 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_8
timestamp 1634918361
transform -1 0 4992 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_9
timestamp 1634918361
transform -1 0 4992 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_10
timestamp 1634918361
transform -1 0 4992 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_11
timestamp 1634918361
transform -1 0 4992 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_12
timestamp 1634918361
transform -1 0 4992 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_13
timestamp 1634918361
transform -1 0 4992 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_14
timestamp 1634918361
transform -1 0 4992 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_15
timestamp 1634918361
transform -1 0 4992 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_16
timestamp 1634918361
transform 1 0 3744 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_17
timestamp 1634918361
transform 1 0 3744 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_18
timestamp 1634918361
transform 1 0 3744 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_19
timestamp 1634918361
transform 1 0 3744 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_20
timestamp 1634918361
transform 1 0 3744 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_21
timestamp 1634918361
transform 1 0 3744 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_22
timestamp 1634918361
transform 1 0 3744 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_23
timestamp 1634918361
transform 1 0 3744 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_24
timestamp 1634918361
transform 1 0 3744 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_25
timestamp 1634918361
transform 1 0 3744 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_26
timestamp 1634918361
transform 1 0 3744 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_27
timestamp 1634918361
transform 1 0 3744 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_28
timestamp 1634918361
transform 1 0 3744 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_29
timestamp 1634918361
transform 1 0 3744 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_30
timestamp 1634918361
transform 1 0 3744 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_31
timestamp 1634918361
transform 1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_32
timestamp 1634918361
transform -1 0 3744 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_33
timestamp 1634918361
transform -1 0 3744 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_34
timestamp 1634918361
transform -1 0 3744 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_35
timestamp 1634918361
transform -1 0 3744 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_36
timestamp 1634918361
transform -1 0 3744 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_37
timestamp 1634918361
transform -1 0 3744 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_38
timestamp 1634918361
transform -1 0 3744 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_39
timestamp 1634918361
transform -1 0 3744 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_40
timestamp 1634918361
transform -1 0 3744 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_41
timestamp 1634918361
transform -1 0 3744 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_42
timestamp 1634918361
transform -1 0 3744 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_43
timestamp 1634918361
transform -1 0 3744 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_44
timestamp 1634918361
transform -1 0 3744 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_45
timestamp 1634918361
transform -1 0 3744 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_46
timestamp 1634918361
transform -1 0 3744 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_47
timestamp 1634918361
transform -1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_48
timestamp 1634918361
transform 1 0 2496 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_49
timestamp 1634918361
transform 1 0 2496 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_50
timestamp 1634918361
transform 1 0 2496 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_51
timestamp 1634918361
transform 1 0 2496 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_52
timestamp 1634918361
transform 1 0 2496 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_53
timestamp 1634918361
transform 1 0 2496 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_54
timestamp 1634918361
transform 1 0 2496 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_55
timestamp 1634918361
transform 1 0 2496 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_56
timestamp 1634918361
transform 1 0 2496 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_57
timestamp 1634918361
transform 1 0 2496 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_58
timestamp 1634918361
transform 1 0 2496 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_59
timestamp 1634918361
transform 1 0 2496 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_60
timestamp 1634918361
transform 1 0 2496 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_61
timestamp 1634918361
transform 1 0 2496 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_62
timestamp 1634918361
transform 1 0 2496 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_63
timestamp 1634918361
transform 1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_64
timestamp 1634918361
transform -1 0 2496 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_65
timestamp 1634918361
transform -1 0 2496 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_66
timestamp 1634918361
transform -1 0 2496 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_67
timestamp 1634918361
transform -1 0 2496 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_68
timestamp 1634918361
transform -1 0 2496 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_69
timestamp 1634918361
transform -1 0 2496 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_70
timestamp 1634918361
transform -1 0 2496 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_71
timestamp 1634918361
transform -1 0 2496 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_72
timestamp 1634918361
transform -1 0 2496 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_73
timestamp 1634918361
transform -1 0 2496 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_74
timestamp 1634918361
transform -1 0 2496 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_75
timestamp 1634918361
transform -1 0 2496 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_76
timestamp 1634918361
transform -1 0 2496 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_77
timestamp 1634918361
transform -1 0 2496 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_78
timestamp 1634918361
transform -1 0 2496 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_79
timestamp 1634918361
transform -1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_80
timestamp 1634918361
transform 1 0 1248 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_81
timestamp 1634918361
transform 1 0 1248 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_82
timestamp 1634918361
transform 1 0 1248 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_83
timestamp 1634918361
transform 1 0 1248 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_84
timestamp 1634918361
transform 1 0 1248 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_85
timestamp 1634918361
transform 1 0 1248 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_86
timestamp 1634918361
transform 1 0 1248 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_87
timestamp 1634918361
transform 1 0 1248 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_88
timestamp 1634918361
transform 1 0 1248 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_89
timestamp 1634918361
transform 1 0 1248 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_90
timestamp 1634918361
transform 1 0 1248 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_91
timestamp 1634918361
transform 1 0 1248 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_92
timestamp 1634918361
transform 1 0 1248 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_93
timestamp 1634918361
transform 1 0 1248 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_94
timestamp 1634918361
transform 1 0 1248 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_95
timestamp 1634918361
transform 1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_96
timestamp 1634918361
transform -1 0 1248 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_97
timestamp 1634918361
transform -1 0 1248 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_98
timestamp 1634918361
transform -1 0 1248 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_99
timestamp 1634918361
transform -1 0 1248 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_100
timestamp 1634918361
transform -1 0 1248 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_101
timestamp 1634918361
transform -1 0 1248 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_102
timestamp 1634918361
transform -1 0 1248 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_103
timestamp 1634918361
transform -1 0 1248 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_104
timestamp 1634918361
transform -1 0 1248 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_105
timestamp 1634918361
transform -1 0 1248 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_106
timestamp 1634918361
transform -1 0 1248 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_107
timestamp 1634918361
transform -1 0 1248 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_108
timestamp 1634918361
transform -1 0 1248 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_109
timestamp 1634918361
transform -1 0 1248 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_110
timestamp 1634918361
transform -1 0 1248 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_111
timestamp 1634918361
transform -1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_112
timestamp 1634918361
transform 1 0 0 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_113
timestamp 1634918361
transform 1 0 0 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_114
timestamp 1634918361
transform 1 0 0 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_115
timestamp 1634918361
transform 1 0 0 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_116
timestamp 1634918361
transform 1 0 0 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_117
timestamp 1634918361
transform 1 0 0 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_118
timestamp 1634918361
transform 1 0 0 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_119
timestamp 1634918361
transform 1 0 0 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_120
timestamp 1634918361
transform 1 0 0 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_121
timestamp 1634918361
transform 1 0 0 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_122
timestamp 1634918361
transform 1 0 0 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_123
timestamp 1634918361
transform 1 0 0 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_124
timestamp 1634918361
transform 1 0 0 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_125
timestamp 1634918361
transform 1 0 0 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_126
timestamp 1634918361
transform 1 0 0 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_127
timestamp 1634918361
transform 1 0 0 0 1 0
box -42 -105 650 421
<< labels >>
rlabel metal1 s 78 0 114 6320 4 bl_0_0
port 1 nsew
rlabel metal1 s 150 0 186 6320 4 br_0_0
port 2 nsew
rlabel metal1 s 294 0 330 6320 4 bl_1_0
port 3 nsew
rlabel metal1 s 366 0 402 6320 4 br_1_0
port 4 nsew
rlabel metal1 s 1134 0 1170 6320 4 bl_0_1
port 5 nsew
rlabel metal1 s 1062 0 1098 6320 4 br_0_1
port 6 nsew
rlabel metal1 s 918 0 954 6320 4 bl_1_1
port 7 nsew
rlabel metal1 s 846 0 882 6320 4 br_1_1
port 8 nsew
rlabel metal1 s 1326 0 1362 6320 4 bl_0_2
port 9 nsew
rlabel metal1 s 1398 0 1434 6320 4 br_0_2
port 10 nsew
rlabel metal1 s 1542 0 1578 6320 4 bl_1_2
port 11 nsew
rlabel metal1 s 1614 0 1650 6320 4 br_1_2
port 12 nsew
rlabel metal1 s 2382 0 2418 6320 4 bl_0_3
port 13 nsew
rlabel metal1 s 2310 0 2346 6320 4 br_0_3
port 14 nsew
rlabel metal1 s 2166 0 2202 6320 4 bl_1_3
port 15 nsew
rlabel metal1 s 2094 0 2130 6320 4 br_1_3
port 16 nsew
rlabel metal1 s 2574 0 2610 6320 4 bl_0_4
port 17 nsew
rlabel metal1 s 2646 0 2682 6320 4 br_0_4
port 18 nsew
rlabel metal1 s 2790 0 2826 6320 4 bl_1_4
port 19 nsew
rlabel metal1 s 2862 0 2898 6320 4 br_1_4
port 20 nsew
rlabel metal1 s 3630 0 3666 6320 4 bl_0_5
port 21 nsew
rlabel metal1 s 3558 0 3594 6320 4 br_0_5
port 22 nsew
rlabel metal1 s 3414 0 3450 6320 4 bl_1_5
port 23 nsew
rlabel metal1 s 3342 0 3378 6320 4 br_1_5
port 24 nsew
rlabel metal1 s 3822 0 3858 6320 4 bl_0_6
port 25 nsew
rlabel metal1 s 3894 0 3930 6320 4 br_0_6
port 26 nsew
rlabel metal1 s 4038 0 4074 6320 4 bl_1_6
port 27 nsew
rlabel metal1 s 4110 0 4146 6320 4 br_1_6
port 28 nsew
rlabel metal1 s 4878 0 4914 6320 4 bl_0_7
port 29 nsew
rlabel metal1 s 4806 0 4842 6320 4 br_0_7
port 30 nsew
rlabel metal1 s 4662 0 4698 6320 4 bl_1_7
port 31 nsew
rlabel metal1 s 4590 0 4626 6320 4 br_1_7
port 32 nsew
rlabel metal2 s 0 323 4992 371 4 wl_0_0
port 33 nsew
rlabel metal2 s 0 103 4992 151 4 wl_1_0
port 34 nsew
rlabel metal2 s 0 419 4992 467 4 wl_0_1
port 35 nsew
rlabel metal2 s 0 639 4992 687 4 wl_1_1
port 36 nsew
rlabel metal2 s 0 1113 4992 1161 4 wl_0_2
port 37 nsew
rlabel metal2 s 0 893 4992 941 4 wl_1_2
port 38 nsew
rlabel metal2 s 0 1209 4992 1257 4 wl_0_3
port 39 nsew
rlabel metal2 s 0 1429 4992 1477 4 wl_1_3
port 40 nsew
rlabel metal2 s 0 1903 4992 1951 4 wl_0_4
port 41 nsew
rlabel metal2 s 0 1683 4992 1731 4 wl_1_4
port 42 nsew
rlabel metal2 s 0 1999 4992 2047 4 wl_0_5
port 43 nsew
rlabel metal2 s 0 2219 4992 2267 4 wl_1_5
port 44 nsew
rlabel metal2 s 0 2693 4992 2741 4 wl_0_6
port 45 nsew
rlabel metal2 s 0 2473 4992 2521 4 wl_1_6
port 46 nsew
rlabel metal2 s 0 2789 4992 2837 4 wl_0_7
port 47 nsew
rlabel metal2 s 0 3009 4992 3057 4 wl_1_7
port 48 nsew
rlabel metal2 s 0 3483 4992 3531 4 wl_0_8
port 49 nsew
rlabel metal2 s 0 3263 4992 3311 4 wl_1_8
port 50 nsew
rlabel metal2 s 0 3579 4992 3627 4 wl_0_9
port 51 nsew
rlabel metal2 s 0 3799 4992 3847 4 wl_1_9
port 52 nsew
rlabel metal2 s 0 4273 4992 4321 4 wl_0_10
port 53 nsew
rlabel metal2 s 0 4053 4992 4101 4 wl_1_10
port 54 nsew
rlabel metal2 s 0 4369 4992 4417 4 wl_0_11
port 55 nsew
rlabel metal2 s 0 4589 4992 4637 4 wl_1_11
port 56 nsew
rlabel metal2 s 0 5063 4992 5111 4 wl_0_12
port 57 nsew
rlabel metal2 s 0 4843 4992 4891 4 wl_1_12
port 58 nsew
rlabel metal2 s 0 5159 4992 5207 4 wl_0_13
port 59 nsew
rlabel metal2 s 0 5379 4992 5427 4 wl_1_13
port 60 nsew
rlabel metal2 s 0 5853 4992 5901 4 wl_0_14
port 61 nsew
rlabel metal2 s 0 5633 4992 5681 4 wl_1_14
port 62 nsew
rlabel metal2 s 0 5949 4992 5997 4 wl_0_15
port 63 nsew
rlabel metal2 s 0 6169 4992 6217 4 wl_1_15
port 64 nsew
rlabel metal1 s 2238 3239 2274 3580 4 vdd
port 65 nsew
rlabel metal1 s 3486 5110 3522 5451 4 vdd
port 65 nsew
rlabel metal1 s 3966 79 4002 420 4 vdd
port 65 nsew
rlabel metal1 s 222 4029 258 4370 4 vdd
port 65 nsew
rlabel metal1 s 3486 79 3522 420 4 vdd
port 65 nsew
rlabel metal1 s 4734 869 4770 1210 4 vdd
port 65 nsew
rlabel metal1 s 2718 3530 2754 3871 4 vdd
port 65 nsew
rlabel metal1 s 2718 3239 2754 3580 4 vdd
port 65 nsew
rlabel metal1 s 2718 1659 2754 2000 4 vdd
port 65 nsew
rlabel metal1 s 3486 1950 3522 2291 4 vdd
port 65 nsew
rlabel metal1 s 2238 5609 2274 5950 4 vdd
port 65 nsew
rlabel metal1 s 3966 3239 4002 3580 4 vdd
port 65 nsew
rlabel metal1 s 3486 5609 3522 5950 4 vdd
port 65 nsew
rlabel metal1 s 2718 4029 2754 4370 4 vdd
port 65 nsew
rlabel metal1 s 2238 1160 2274 1501 4 vdd
port 65 nsew
rlabel metal1 s 3486 2449 3522 2790 4 vdd
port 65 nsew
rlabel metal1 s 2718 1950 2754 2291 4 vdd
port 65 nsew
rlabel metal1 s 990 370 1026 711 4 vdd
port 65 nsew
rlabel metal1 s 3966 5110 4002 5451 4 vdd
port 65 nsew
rlabel metal1 s 3486 3530 3522 3871 4 vdd
port 65 nsew
rlabel metal1 s 2718 2740 2754 3081 4 vdd
port 65 nsew
rlabel metal1 s 3966 1160 4002 1501 4 vdd
port 65 nsew
rlabel metal1 s 3966 1950 4002 2291 4 vdd
port 65 nsew
rlabel metal1 s 3486 4819 3522 5160 4 vdd
port 65 nsew
rlabel metal1 s 990 3239 1026 3580 4 vdd
port 65 nsew
rlabel metal1 s 990 1950 1026 2291 4 vdd
port 65 nsew
rlabel metal1 s 4734 2740 4770 3081 4 vdd
port 65 nsew
rlabel metal1 s 3486 2740 3522 3081 4 vdd
port 65 nsew
rlabel metal1 s 2718 5900 2754 6241 4 vdd
port 65 nsew
rlabel metal1 s 1470 5110 1506 5451 4 vdd
port 65 nsew
rlabel metal1 s 4734 4819 4770 5160 4 vdd
port 65 nsew
rlabel metal1 s 1470 3530 1506 3871 4 vdd
port 65 nsew
rlabel metal1 s 1470 5609 1506 5950 4 vdd
port 65 nsew
rlabel metal1 s 2718 1160 2754 1501 4 vdd
port 65 nsew
rlabel metal1 s 3966 2740 4002 3081 4 vdd
port 65 nsew
rlabel metal1 s 1470 4320 1506 4661 4 vdd
port 65 nsew
rlabel metal1 s 2238 4320 2274 4661 4 vdd
port 65 nsew
rlabel metal1 s 3966 4819 4002 5160 4 vdd
port 65 nsew
rlabel metal1 s 222 1659 258 2000 4 vdd
port 65 nsew
rlabel metal1 s 3966 2449 4002 2790 4 vdd
port 65 nsew
rlabel metal1 s 4734 4029 4770 4370 4 vdd
port 65 nsew
rlabel metal1 s 1470 1160 1506 1501 4 vdd
port 65 nsew
rlabel metal1 s 3486 1659 3522 2000 4 vdd
port 65 nsew
rlabel metal1 s 4734 79 4770 420 4 vdd
port 65 nsew
rlabel metal1 s 990 4320 1026 4661 4 vdd
port 65 nsew
rlabel metal1 s 2718 2449 2754 2790 4 vdd
port 65 nsew
rlabel metal1 s 1470 1950 1506 2291 4 vdd
port 65 nsew
rlabel metal1 s 990 5609 1026 5950 4 vdd
port 65 nsew
rlabel metal1 s 3966 5900 4002 6241 4 vdd
port 65 nsew
rlabel metal1 s 3966 1659 4002 2000 4 vdd
port 65 nsew
rlabel metal1 s 990 79 1026 420 4 vdd
port 65 nsew
rlabel metal1 s 990 2740 1026 3081 4 vdd
port 65 nsew
rlabel metal1 s 990 2449 1026 2790 4 vdd
port 65 nsew
rlabel metal1 s 4734 5900 4770 6241 4 vdd
port 65 nsew
rlabel metal1 s 3966 370 4002 711 4 vdd
port 65 nsew
rlabel metal1 s 2718 4819 2754 5160 4 vdd
port 65 nsew
rlabel metal1 s 4734 5609 4770 5950 4 vdd
port 65 nsew
rlabel metal1 s 3486 4320 3522 4661 4 vdd
port 65 nsew
rlabel metal1 s 222 4819 258 5160 4 vdd
port 65 nsew
rlabel metal1 s 2238 869 2274 1210 4 vdd
port 65 nsew
rlabel metal1 s 3966 4320 4002 4661 4 vdd
port 65 nsew
rlabel metal1 s 3966 3530 4002 3871 4 vdd
port 65 nsew
rlabel metal1 s 1470 4819 1506 5160 4 vdd
port 65 nsew
rlabel metal1 s 2238 79 2274 420 4 vdd
port 65 nsew
rlabel metal1 s 990 5900 1026 6241 4 vdd
port 65 nsew
rlabel metal1 s 222 370 258 711 4 vdd
port 65 nsew
rlabel metal1 s 2238 5900 2274 6241 4 vdd
port 65 nsew
rlabel metal1 s 4734 3530 4770 3871 4 vdd
port 65 nsew
rlabel metal1 s 222 2740 258 3081 4 vdd
port 65 nsew
rlabel metal1 s 4734 1160 4770 1501 4 vdd
port 65 nsew
rlabel metal1 s 3486 370 3522 711 4 vdd
port 65 nsew
rlabel metal1 s 2718 869 2754 1210 4 vdd
port 65 nsew
rlabel metal1 s 222 1160 258 1501 4 vdd
port 65 nsew
rlabel metal1 s 2238 370 2274 711 4 vdd
port 65 nsew
rlabel metal1 s 2718 5110 2754 5451 4 vdd
port 65 nsew
rlabel metal1 s 2718 4320 2754 4661 4 vdd
port 65 nsew
rlabel metal1 s 2238 3530 2274 3871 4 vdd
port 65 nsew
rlabel metal1 s 990 3530 1026 3871 4 vdd
port 65 nsew
rlabel metal1 s 1470 3239 1506 3580 4 vdd
port 65 nsew
rlabel metal1 s 2718 370 2754 711 4 vdd
port 65 nsew
rlabel metal1 s 222 5110 258 5451 4 vdd
port 65 nsew
rlabel metal1 s 1470 2740 1506 3081 4 vdd
port 65 nsew
rlabel metal1 s 2238 4029 2274 4370 4 vdd
port 65 nsew
rlabel metal1 s 4734 1659 4770 2000 4 vdd
port 65 nsew
rlabel metal1 s 2238 1950 2274 2291 4 vdd
port 65 nsew
rlabel metal1 s 3486 869 3522 1210 4 vdd
port 65 nsew
rlabel metal1 s 1470 79 1506 420 4 vdd
port 65 nsew
rlabel metal1 s 3966 4029 4002 4370 4 vdd
port 65 nsew
rlabel metal1 s 222 1950 258 2291 4 vdd
port 65 nsew
rlabel metal1 s 1470 370 1506 711 4 vdd
port 65 nsew
rlabel metal1 s 1470 2449 1506 2790 4 vdd
port 65 nsew
rlabel metal1 s 2238 1659 2274 2000 4 vdd
port 65 nsew
rlabel metal1 s 2238 2449 2274 2790 4 vdd
port 65 nsew
rlabel metal1 s 4734 3239 4770 3580 4 vdd
port 65 nsew
rlabel metal1 s 222 3530 258 3871 4 vdd
port 65 nsew
rlabel metal1 s 4734 5110 4770 5451 4 vdd
port 65 nsew
rlabel metal1 s 222 5900 258 6241 4 vdd
port 65 nsew
rlabel metal1 s 4734 370 4770 711 4 vdd
port 65 nsew
rlabel metal1 s 4734 4320 4770 4661 4 vdd
port 65 nsew
rlabel metal1 s 222 5609 258 5950 4 vdd
port 65 nsew
rlabel metal1 s 990 4819 1026 5160 4 vdd
port 65 nsew
rlabel metal1 s 990 1160 1026 1501 4 vdd
port 65 nsew
rlabel metal1 s 2238 4819 2274 5160 4 vdd
port 65 nsew
rlabel metal1 s 2718 79 2754 420 4 vdd
port 65 nsew
rlabel metal1 s 990 4029 1026 4370 4 vdd
port 65 nsew
rlabel metal1 s 990 5110 1026 5451 4 vdd
port 65 nsew
rlabel metal1 s 222 79 258 420 4 vdd
port 65 nsew
rlabel metal1 s 2238 2740 2274 3081 4 vdd
port 65 nsew
rlabel metal1 s 990 869 1026 1210 4 vdd
port 65 nsew
rlabel metal1 s 4734 2449 4770 2790 4 vdd
port 65 nsew
rlabel metal1 s 1470 4029 1506 4370 4 vdd
port 65 nsew
rlabel metal1 s 3966 869 4002 1210 4 vdd
port 65 nsew
rlabel metal1 s 1470 869 1506 1210 4 vdd
port 65 nsew
rlabel metal1 s 222 4320 258 4661 4 vdd
port 65 nsew
rlabel metal1 s 222 3239 258 3580 4 vdd
port 65 nsew
rlabel metal1 s 222 869 258 1210 4 vdd
port 65 nsew
rlabel metal1 s 222 2449 258 2790 4 vdd
port 65 nsew
rlabel metal1 s 3486 4029 3522 4370 4 vdd
port 65 nsew
rlabel metal1 s 2238 5110 2274 5451 4 vdd
port 65 nsew
rlabel metal1 s 1470 5900 1506 6241 4 vdd
port 65 nsew
rlabel metal1 s 2718 5609 2754 5950 4 vdd
port 65 nsew
rlabel metal1 s 1470 1659 1506 2000 4 vdd
port 65 nsew
rlabel metal1 s 4734 1950 4770 2291 4 vdd
port 65 nsew
rlabel metal1 s 3966 5609 4002 5950 4 vdd
port 65 nsew
rlabel metal1 s 3486 1160 3522 1501 4 vdd
port 65 nsew
rlabel metal1 s 3486 5900 3522 6241 4 vdd
port 65 nsew
rlabel metal1 s 3486 3239 3522 3580 4 vdd
port 65 nsew
rlabel metal1 s 990 1659 1026 2000 4 vdd
port 65 nsew
rlabel metal2 s 2682 -55 2790 55 4 gnd
port 66 nsew
rlabel metal2 s 4698 2095 4806 2171 4 gnd
port 66 nsew
rlabel metal2 s 3930 199 4038 275 4 gnd
port 66 nsew
rlabel metal2 s 3450 2095 3558 2171 4 gnd
port 66 nsew
rlabel metal2 s 3450 1779 3558 1855 4 gnd
port 66 nsew
rlabel metal2 s 3450 735 3558 845 4 gnd
port 66 nsew
rlabel metal2 s 4698 4685 4806 4795 4 gnd
port 66 nsew
rlabel metal2 s 186 1525 294 1635 4 gnd
port 66 nsew
rlabel metal2 s 3450 2885 3558 2961 4 gnd
port 66 nsew
rlabel metal2 s 3930 3675 4038 3751 4 gnd
port 66 nsew
rlabel metal2 s 186 4149 294 4225 4 gnd
port 66 nsew
rlabel metal2 s 4698 4939 4806 5015 4 gnd
port 66 nsew
rlabel metal2 s 1434 5729 1542 5805 4 gnd
port 66 nsew
rlabel metal2 s 4698 6265 4806 6375 4 gnd
port 66 nsew
rlabel metal2 s 4698 2315 4806 2425 4 gnd
port 66 nsew
rlabel metal2 s 186 1305 294 1381 4 gnd
port 66 nsew
rlabel metal2 s 3450 1525 3558 1635 4 gnd
port 66 nsew
rlabel metal2 s 4698 1779 4806 1855 4 gnd
port 66 nsew
rlabel metal2 s 2202 2095 2310 2171 4 gnd
port 66 nsew
rlabel metal2 s 4698 2885 4806 2961 4 gnd
port 66 nsew
rlabel metal2 s 3450 3895 3558 4005 4 gnd
port 66 nsew
rlabel metal2 s 3930 3895 4038 4005 4 gnd
port 66 nsew
rlabel metal2 s 3930 4939 4038 5015 4 gnd
port 66 nsew
rlabel metal2 s 2202 5255 2310 5331 4 gnd
port 66 nsew
rlabel metal2 s 3930 5475 4038 5585 4 gnd
port 66 nsew
rlabel metal2 s 2202 3895 2310 4005 4 gnd
port 66 nsew
rlabel metal2 s 2202 4149 2310 4225 4 gnd
port 66 nsew
rlabel metal2 s 186 1779 294 1855 4 gnd
port 66 nsew
rlabel metal2 s 954 5475 1062 5585 4 gnd
port 66 nsew
rlabel metal2 s 2202 5475 2310 5585 4 gnd
port 66 nsew
rlabel metal2 s 2682 1779 2790 1855 4 gnd
port 66 nsew
rlabel metal2 s 954 3359 1062 3435 4 gnd
port 66 nsew
rlabel metal2 s 3930 1305 4038 1381 4 gnd
port 66 nsew
rlabel metal2 s 2202 735 2310 845 4 gnd
port 66 nsew
rlabel metal2 s 3450 989 3558 1065 4 gnd
port 66 nsew
rlabel metal2 s 2682 4149 2790 4225 4 gnd
port 66 nsew
rlabel metal2 s 186 5475 294 5585 4 gnd
port 66 nsew
rlabel metal2 s 954 4149 1062 4225 4 gnd
port 66 nsew
rlabel metal2 s 1434 5475 1542 5585 4 gnd
port 66 nsew
rlabel metal2 s 954 2885 1062 2961 4 gnd
port 66 nsew
rlabel metal2 s 3930 6265 4038 6375 4 gnd
port 66 nsew
rlabel metal2 s 4698 989 4806 1065 4 gnd
port 66 nsew
rlabel metal2 s 2682 3105 2790 3215 4 gnd
port 66 nsew
rlabel metal2 s 3930 3105 4038 3215 4 gnd
port 66 nsew
rlabel metal2 s 1434 2885 1542 2961 4 gnd
port 66 nsew
rlabel metal2 s 4698 1305 4806 1381 4 gnd
port 66 nsew
rlabel metal2 s 186 199 294 275 4 gnd
port 66 nsew
rlabel metal2 s 186 989 294 1065 4 gnd
port 66 nsew
rlabel metal2 s 186 4939 294 5015 4 gnd
port 66 nsew
rlabel metal2 s 2682 5729 2790 5805 4 gnd
port 66 nsew
rlabel metal2 s 954 6045 1062 6121 4 gnd
port 66 nsew
rlabel metal2 s 2682 4465 2790 4541 4 gnd
port 66 nsew
rlabel metal2 s 1434 1779 1542 1855 4 gnd
port 66 nsew
rlabel metal2 s 186 2569 294 2645 4 gnd
port 66 nsew
rlabel metal2 s 2202 4685 2310 4795 4 gnd
port 66 nsew
rlabel metal2 s 4698 5255 4806 5331 4 gnd
port 66 nsew
rlabel metal2 s 1434 4465 1542 4541 4 gnd
port 66 nsew
rlabel metal2 s 1434 1525 1542 1635 4 gnd
port 66 nsew
rlabel metal2 s 186 -55 294 55 4 gnd
port 66 nsew
rlabel metal2 s 3930 989 4038 1065 4 gnd
port 66 nsew
rlabel metal2 s 954 5729 1062 5805 4 gnd
port 66 nsew
rlabel metal2 s 4698 1525 4806 1635 4 gnd
port 66 nsew
rlabel metal2 s 3450 4465 3558 4541 4 gnd
port 66 nsew
rlabel metal2 s 954 1305 1062 1381 4 gnd
port 66 nsew
rlabel metal2 s 2202 515 2310 591 4 gnd
port 66 nsew
rlabel metal2 s 3930 4465 4038 4541 4 gnd
port 66 nsew
rlabel metal2 s 2202 1305 2310 1381 4 gnd
port 66 nsew
rlabel metal2 s 186 515 294 591 4 gnd
port 66 nsew
rlabel metal2 s 2202 2885 2310 2961 4 gnd
port 66 nsew
rlabel metal2 s 3450 5729 3558 5805 4 gnd
port 66 nsew
rlabel metal2 s 3930 1779 4038 1855 4 gnd
port 66 nsew
rlabel metal2 s 954 4465 1062 4541 4 gnd
port 66 nsew
rlabel metal2 s 186 6265 294 6375 4 gnd
port 66 nsew
rlabel metal2 s 1434 735 1542 845 4 gnd
port 66 nsew
rlabel metal2 s 954 1525 1062 1635 4 gnd
port 66 nsew
rlabel metal2 s 2682 735 2790 845 4 gnd
port 66 nsew
rlabel metal2 s 186 3895 294 4005 4 gnd
port 66 nsew
rlabel metal2 s 1434 5255 1542 5331 4 gnd
port 66 nsew
rlabel metal2 s 2202 989 2310 1065 4 gnd
port 66 nsew
rlabel metal2 s 954 735 1062 845 4 gnd
port 66 nsew
rlabel metal2 s 186 6045 294 6121 4 gnd
port 66 nsew
rlabel metal2 s 2202 2315 2310 2425 4 gnd
port 66 nsew
rlabel metal2 s 3930 2885 4038 2961 4 gnd
port 66 nsew
rlabel metal2 s 3450 2315 3558 2425 4 gnd
port 66 nsew
rlabel metal2 s 3450 -55 3558 55 4 gnd
port 66 nsew
rlabel metal2 s 2682 3895 2790 4005 4 gnd
port 66 nsew
rlabel metal2 s 186 3105 294 3215 4 gnd
port 66 nsew
rlabel metal2 s 3450 6265 3558 6375 4 gnd
port 66 nsew
rlabel metal2 s 4698 3359 4806 3435 4 gnd
port 66 nsew
rlabel metal2 s 2682 4939 2790 5015 4 gnd
port 66 nsew
rlabel metal2 s 2202 4939 2310 5015 4 gnd
port 66 nsew
rlabel metal2 s 186 2315 294 2425 4 gnd
port 66 nsew
rlabel metal2 s 1434 4939 1542 5015 4 gnd
port 66 nsew
rlabel metal2 s 4698 735 4806 845 4 gnd
port 66 nsew
rlabel metal2 s 4698 -55 4806 55 4 gnd
port 66 nsew
rlabel metal2 s 3930 5729 4038 5805 4 gnd
port 66 nsew
rlabel metal2 s 3930 2569 4038 2645 4 gnd
port 66 nsew
rlabel metal2 s 2682 6265 2790 6375 4 gnd
port 66 nsew
rlabel metal2 s 954 989 1062 1065 4 gnd
port 66 nsew
rlabel metal2 s 3930 3359 4038 3435 4 gnd
port 66 nsew
rlabel metal2 s 186 5255 294 5331 4 gnd
port 66 nsew
rlabel metal2 s 954 4685 1062 4795 4 gnd
port 66 nsew
rlabel metal2 s 186 3675 294 3751 4 gnd
port 66 nsew
rlabel metal2 s 1434 515 1542 591 4 gnd
port 66 nsew
rlabel metal2 s 2682 5255 2790 5331 4 gnd
port 66 nsew
rlabel metal2 s 1434 6045 1542 6121 4 gnd
port 66 nsew
rlabel metal2 s 3930 2315 4038 2425 4 gnd
port 66 nsew
rlabel metal2 s 2202 3105 2310 3215 4 gnd
port 66 nsew
rlabel metal2 s 954 6265 1062 6375 4 gnd
port 66 nsew
rlabel metal2 s 954 2095 1062 2171 4 gnd
port 66 nsew
rlabel metal2 s 4698 5729 4806 5805 4 gnd
port 66 nsew
rlabel metal2 s 2682 5475 2790 5585 4 gnd
port 66 nsew
rlabel metal2 s 4698 6045 4806 6121 4 gnd
port 66 nsew
rlabel metal2 s 2682 2095 2790 2171 4 gnd
port 66 nsew
rlabel metal2 s 3930 2095 4038 2171 4 gnd
port 66 nsew
rlabel metal2 s 3930 -55 4038 55 4 gnd
port 66 nsew
rlabel metal2 s 954 515 1062 591 4 gnd
port 66 nsew
rlabel metal2 s 4698 3105 4806 3215 4 gnd
port 66 nsew
rlabel metal2 s 3930 4149 4038 4225 4 gnd
port 66 nsew
rlabel metal2 s 1434 2095 1542 2171 4 gnd
port 66 nsew
rlabel metal2 s 954 3895 1062 4005 4 gnd
port 66 nsew
rlabel metal2 s 3930 515 4038 591 4 gnd
port 66 nsew
rlabel metal2 s 3450 1305 3558 1381 4 gnd
port 66 nsew
rlabel metal2 s 1434 3895 1542 4005 4 gnd
port 66 nsew
rlabel metal2 s 186 3359 294 3435 4 gnd
port 66 nsew
rlabel metal2 s 1434 6265 1542 6375 4 gnd
port 66 nsew
rlabel metal2 s 2202 6045 2310 6121 4 gnd
port 66 nsew
rlabel metal2 s 2682 3359 2790 3435 4 gnd
port 66 nsew
rlabel metal2 s 4698 4149 4806 4225 4 gnd
port 66 nsew
rlabel metal2 s 3450 199 3558 275 4 gnd
port 66 nsew
rlabel metal2 s 186 735 294 845 4 gnd
port 66 nsew
rlabel metal2 s 2682 2885 2790 2961 4 gnd
port 66 nsew
rlabel metal2 s 3450 4149 3558 4225 4 gnd
port 66 nsew
rlabel metal2 s 954 3675 1062 3751 4 gnd
port 66 nsew
rlabel metal2 s 3930 5255 4038 5331 4 gnd
port 66 nsew
rlabel metal2 s 4698 2569 4806 2645 4 gnd
port 66 nsew
rlabel metal2 s 2682 2569 2790 2645 4 gnd
port 66 nsew
rlabel metal2 s 3450 4685 3558 4795 4 gnd
port 66 nsew
rlabel metal2 s 4698 3675 4806 3751 4 gnd
port 66 nsew
rlabel metal2 s 3930 735 4038 845 4 gnd
port 66 nsew
rlabel metal2 s 2202 1525 2310 1635 4 gnd
port 66 nsew
rlabel metal2 s 2682 199 2790 275 4 gnd
port 66 nsew
rlabel metal2 s 1434 2569 1542 2645 4 gnd
port 66 nsew
rlabel metal2 s 4698 3895 4806 4005 4 gnd
port 66 nsew
rlabel metal2 s 3450 5255 3558 5331 4 gnd
port 66 nsew
rlabel metal2 s 3450 4939 3558 5015 4 gnd
port 66 nsew
rlabel metal2 s 3450 515 3558 591 4 gnd
port 66 nsew
rlabel metal2 s 186 5729 294 5805 4 gnd
port 66 nsew
rlabel metal2 s 3930 1525 4038 1635 4 gnd
port 66 nsew
rlabel metal2 s 1434 2315 1542 2425 4 gnd
port 66 nsew
rlabel metal2 s 186 2885 294 2961 4 gnd
port 66 nsew
rlabel metal2 s 3450 3675 3558 3751 4 gnd
port 66 nsew
rlabel metal2 s 4698 4465 4806 4541 4 gnd
port 66 nsew
rlabel metal2 s 2682 6045 2790 6121 4 gnd
port 66 nsew
rlabel metal2 s 2202 6265 2310 6375 4 gnd
port 66 nsew
rlabel metal2 s 3450 2569 3558 2645 4 gnd
port 66 nsew
rlabel metal2 s 2682 989 2790 1065 4 gnd
port 66 nsew
rlabel metal2 s 3450 3359 3558 3435 4 gnd
port 66 nsew
rlabel metal2 s 2682 1305 2790 1381 4 gnd
port 66 nsew
rlabel metal2 s 2682 3675 2790 3751 4 gnd
port 66 nsew
rlabel metal2 s 2682 1525 2790 1635 4 gnd
port 66 nsew
rlabel metal2 s 2202 3675 2310 3751 4 gnd
port 66 nsew
rlabel metal2 s 4698 199 4806 275 4 gnd
port 66 nsew
rlabel metal2 s 954 1779 1062 1855 4 gnd
port 66 nsew
rlabel metal2 s 954 4939 1062 5015 4 gnd
port 66 nsew
rlabel metal2 s 186 4685 294 4795 4 gnd
port 66 nsew
rlabel metal2 s 1434 4685 1542 4795 4 gnd
port 66 nsew
rlabel metal2 s 2202 1779 2310 1855 4 gnd
port 66 nsew
rlabel metal2 s 954 2569 1062 2645 4 gnd
port 66 nsew
rlabel metal2 s 2202 2569 2310 2645 4 gnd
port 66 nsew
rlabel metal2 s 2202 3359 2310 3435 4 gnd
port 66 nsew
rlabel metal2 s 1434 4149 1542 4225 4 gnd
port 66 nsew
rlabel metal2 s 2202 199 2310 275 4 gnd
port 66 nsew
rlabel metal2 s 1434 3105 1542 3215 4 gnd
port 66 nsew
rlabel metal2 s 4698 515 4806 591 4 gnd
port 66 nsew
rlabel metal2 s 3450 6045 3558 6121 4 gnd
port 66 nsew
rlabel metal2 s 1434 989 1542 1065 4 gnd
port 66 nsew
rlabel metal2 s 2202 5729 2310 5805 4 gnd
port 66 nsew
rlabel metal2 s 2202 4465 2310 4541 4 gnd
port 66 nsew
rlabel metal2 s 3930 6045 4038 6121 4 gnd
port 66 nsew
rlabel metal2 s 1434 1305 1542 1381 4 gnd
port 66 nsew
rlabel metal2 s 1434 199 1542 275 4 gnd
port 66 nsew
rlabel metal2 s 954 199 1062 275 4 gnd
port 66 nsew
rlabel metal2 s 1434 3675 1542 3751 4 gnd
port 66 nsew
rlabel metal2 s 3930 4685 4038 4795 4 gnd
port 66 nsew
rlabel metal2 s 2682 4685 2790 4795 4 gnd
port 66 nsew
rlabel metal2 s 954 5255 1062 5331 4 gnd
port 66 nsew
rlabel metal2 s 186 2095 294 2171 4 gnd
port 66 nsew
rlabel metal2 s 1434 3359 1542 3435 4 gnd
port 66 nsew
rlabel metal2 s 3450 3105 3558 3215 4 gnd
port 66 nsew
rlabel metal2 s 186 4465 294 4541 4 gnd
port 66 nsew
rlabel metal2 s 4698 5475 4806 5585 4 gnd
port 66 nsew
rlabel metal2 s 1434 -55 1542 55 4 gnd
port 66 nsew
rlabel metal2 s 954 3105 1062 3215 4 gnd
port 66 nsew
rlabel metal2 s 3450 5475 3558 5585 4 gnd
port 66 nsew
rlabel metal2 s 954 -55 1062 55 4 gnd
port 66 nsew
rlabel metal2 s 2202 -55 2310 55 4 gnd
port 66 nsew
rlabel metal2 s 2682 515 2790 591 4 gnd
port 66 nsew
rlabel metal2 s 2682 2315 2790 2425 4 gnd
port 66 nsew
rlabel metal2 s 954 2315 1062 2425 4 gnd
port 66 nsew
<< properties >>
string FIXED_BBOX 0 0 4992 6320
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 582702
string GDS_START 505250
<< end >>
