magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1296 -1309 10640 2727
<< locali >>
rect 567 1431 601 1447
rect 567 1381 601 1397
rect 1735 1431 1769 1447
rect 1735 1381 1769 1397
rect 2903 1431 2937 1447
rect 2903 1381 2937 1397
rect 4071 1431 4105 1447
rect 4071 1381 4105 1397
rect 5239 1431 5273 1447
rect 5239 1381 5273 1397
rect 6407 1431 6441 1447
rect 6407 1381 6441 1397
rect 7575 1431 7609 1447
rect 7575 1381 7609 1397
rect 8743 1431 8777 1447
rect 8743 1381 8777 1397
rect 567 17 601 33
rect 567 -33 601 -17
rect 1735 17 1769 33
rect 1735 -33 1769 -17
rect 2903 17 2937 33
rect 2903 -33 2937 -17
rect 4071 17 4105 33
rect 4071 -33 4105 -17
rect 5239 17 5273 33
rect 5239 -33 5273 -17
rect 6407 17 6441 33
rect 6407 -33 6441 -17
rect 7575 17 7609 33
rect 7575 -33 7609 -17
rect 8743 17 8777 33
rect 8743 -33 8777 -17
<< viali >>
rect 567 1397 601 1431
rect 1735 1397 1769 1431
rect 2903 1397 2937 1431
rect 4071 1397 4105 1431
rect 5239 1397 5273 1431
rect 6407 1397 6441 1431
rect 7575 1397 7609 1431
rect 8743 1397 8777 1431
rect 567 -17 601 17
rect 1735 -17 1769 17
rect 2903 -17 2937 17
rect 4071 -17 4105 17
rect 5239 -17 5273 17
rect 6407 -17 6441 17
rect 7575 -17 7609 17
rect 8743 -17 8777 17
<< metal1 >>
rect 552 1388 558 1440
rect 610 1388 616 1440
rect 1720 1388 1726 1440
rect 1778 1388 1784 1440
rect 2888 1388 2894 1440
rect 2946 1388 2952 1440
rect 4056 1388 4062 1440
rect 4114 1388 4120 1440
rect 5224 1388 5230 1440
rect 5282 1388 5288 1440
rect 6392 1388 6398 1440
rect 6450 1388 6456 1440
rect 7560 1388 7566 1440
rect 7618 1388 7624 1440
rect 8728 1388 8734 1440
rect 8786 1388 8792 1440
rect 552 -26 558 26
rect 610 -26 616 26
rect 1720 -26 1726 26
rect 1778 -26 1784 26
rect 2888 -26 2894 26
rect 2946 -26 2952 26
rect 4056 -26 4062 26
rect 4114 -26 4120 26
rect 5224 -26 5230 26
rect 5282 -26 5288 26
rect 6392 -26 6398 26
rect 6450 -26 6456 26
rect 7560 -26 7566 26
rect 7618 -26 7624 26
rect 8728 -26 8734 26
rect 8786 -26 8792 26
<< via1 >>
rect 558 1431 610 1440
rect 558 1397 567 1431
rect 567 1397 601 1431
rect 601 1397 610 1431
rect 558 1388 610 1397
rect 1726 1431 1778 1440
rect 1726 1397 1735 1431
rect 1735 1397 1769 1431
rect 1769 1397 1778 1431
rect 1726 1388 1778 1397
rect 2894 1431 2946 1440
rect 2894 1397 2903 1431
rect 2903 1397 2937 1431
rect 2937 1397 2946 1431
rect 2894 1388 2946 1397
rect 4062 1431 4114 1440
rect 4062 1397 4071 1431
rect 4071 1397 4105 1431
rect 4105 1397 4114 1431
rect 4062 1388 4114 1397
rect 5230 1431 5282 1440
rect 5230 1397 5239 1431
rect 5239 1397 5273 1431
rect 5273 1397 5282 1431
rect 5230 1388 5282 1397
rect 6398 1431 6450 1440
rect 6398 1397 6407 1431
rect 6407 1397 6441 1431
rect 6441 1397 6450 1431
rect 6398 1388 6450 1397
rect 7566 1431 7618 1440
rect 7566 1397 7575 1431
rect 7575 1397 7609 1431
rect 7609 1397 7618 1431
rect 7566 1388 7618 1397
rect 8734 1431 8786 1440
rect 8734 1397 8743 1431
rect 8743 1397 8777 1431
rect 8777 1397 8786 1431
rect 8734 1388 8786 1397
rect 558 17 610 26
rect 558 -17 567 17
rect 567 -17 601 17
rect 601 -17 610 17
rect 558 -26 610 -17
rect 1726 17 1778 26
rect 1726 -17 1735 17
rect 1735 -17 1769 17
rect 1769 -17 1778 17
rect 1726 -26 1778 -17
rect 2894 17 2946 26
rect 2894 -17 2903 17
rect 2903 -17 2937 17
rect 2937 -17 2946 17
rect 2894 -26 2946 -17
rect 4062 17 4114 26
rect 4062 -17 4071 17
rect 4071 -17 4105 17
rect 4105 -17 4114 17
rect 4062 -26 4114 -17
rect 5230 17 5282 26
rect 5230 -17 5239 17
rect 5239 -17 5273 17
rect 5273 -17 5282 17
rect 5230 -26 5282 -17
rect 6398 17 6450 26
rect 6398 -17 6407 17
rect 6407 -17 6441 17
rect 6441 -17 6450 17
rect 6398 -26 6450 -17
rect 7566 17 7618 26
rect 7566 -17 7575 17
rect 7575 -17 7609 17
rect 7609 -17 7618 17
rect 7566 -26 7618 -17
rect 8734 17 8786 26
rect 8734 -17 8743 17
rect 8743 -17 8777 17
rect 8777 -17 8786 17
rect 8734 -26 8786 -17
<< metal2 >>
rect 556 1442 612 1451
rect 137 538 203 590
rect 369 345 397 1414
rect 1724 1442 1780 1451
rect 556 1377 612 1386
rect 1082 609 1148 661
rect 1305 538 1371 590
rect 1537 345 1565 1414
rect 2892 1442 2948 1451
rect 1724 1377 1780 1386
rect 2250 609 2316 661
rect 2473 538 2539 590
rect 2705 345 2733 1414
rect 4060 1442 4116 1451
rect 2892 1377 2948 1386
rect 3418 609 3484 661
rect 3641 538 3707 590
rect 3873 345 3901 1414
rect 5228 1442 5284 1451
rect 4060 1377 4116 1386
rect 4586 609 4652 661
rect 4809 538 4875 590
rect 5041 345 5069 1414
rect 6396 1442 6452 1451
rect 5228 1377 5284 1386
rect 5754 609 5820 661
rect 5977 538 6043 590
rect 6209 345 6237 1414
rect 7564 1442 7620 1451
rect 6396 1377 6452 1386
rect 6922 609 6988 661
rect 7145 538 7211 590
rect 7377 345 7405 1414
rect 8732 1442 8788 1451
rect 7564 1377 7620 1386
rect 8090 609 8156 661
rect 8313 538 8379 590
rect 8545 345 8573 1414
rect 8732 1377 8788 1386
rect 9258 609 9324 661
rect 368 336 424 345
rect 368 271 424 280
rect 1536 336 1592 345
rect 1536 271 1592 280
rect 2704 336 2760 345
rect 2704 271 2760 280
rect 3872 336 3928 345
rect 3872 271 3928 280
rect 5040 336 5096 345
rect 5040 271 5096 280
rect 6208 336 6264 345
rect 6208 271 6264 280
rect 7376 336 7432 345
rect 7376 271 7432 280
rect 8544 336 8600 345
rect 8544 271 8600 280
rect 369 0 397 271
rect 556 28 612 37
rect 1537 0 1565 271
rect 1724 28 1780 37
rect 556 -37 612 -28
rect 2705 0 2733 271
rect 2892 28 2948 37
rect 1724 -37 1780 -28
rect 3873 0 3901 271
rect 4060 28 4116 37
rect 2892 -37 2948 -28
rect 5041 0 5069 271
rect 5228 28 5284 37
rect 4060 -37 4116 -28
rect 6209 0 6237 271
rect 6396 28 6452 37
rect 5228 -37 5284 -28
rect 7377 0 7405 271
rect 7564 28 7620 37
rect 6396 -37 6452 -28
rect 8545 0 8573 271
rect 8732 28 8788 37
rect 7564 -37 7620 -28
rect 8732 -37 8788 -28
<< via2 >>
rect 556 1440 612 1442
rect 556 1388 558 1440
rect 558 1388 610 1440
rect 610 1388 612 1440
rect 1724 1440 1780 1442
rect 556 1386 612 1388
rect 1724 1388 1726 1440
rect 1726 1388 1778 1440
rect 1778 1388 1780 1440
rect 2892 1440 2948 1442
rect 1724 1386 1780 1388
rect 2892 1388 2894 1440
rect 2894 1388 2946 1440
rect 2946 1388 2948 1440
rect 4060 1440 4116 1442
rect 2892 1386 2948 1388
rect 4060 1388 4062 1440
rect 4062 1388 4114 1440
rect 4114 1388 4116 1440
rect 5228 1440 5284 1442
rect 4060 1386 4116 1388
rect 5228 1388 5230 1440
rect 5230 1388 5282 1440
rect 5282 1388 5284 1440
rect 6396 1440 6452 1442
rect 5228 1386 5284 1388
rect 6396 1388 6398 1440
rect 6398 1388 6450 1440
rect 6450 1388 6452 1440
rect 7564 1440 7620 1442
rect 6396 1386 6452 1388
rect 7564 1388 7566 1440
rect 7566 1388 7618 1440
rect 7618 1388 7620 1440
rect 8732 1440 8788 1442
rect 7564 1386 7620 1388
rect 8732 1388 8734 1440
rect 8734 1388 8786 1440
rect 8786 1388 8788 1440
rect 8732 1386 8788 1388
rect 368 280 424 336
rect 1536 280 1592 336
rect 2704 280 2760 336
rect 3872 280 3928 336
rect 5040 280 5096 336
rect 6208 280 6264 336
rect 7376 280 7432 336
rect 8544 280 8600 336
rect 556 26 612 28
rect 556 -26 558 26
rect 558 -26 610 26
rect 610 -26 612 26
rect 1724 26 1780 28
rect 556 -28 612 -26
rect 1724 -26 1726 26
rect 1726 -26 1778 26
rect 1778 -26 1780 26
rect 2892 26 2948 28
rect 1724 -28 1780 -26
rect 2892 -26 2894 26
rect 2894 -26 2946 26
rect 2946 -26 2948 26
rect 4060 26 4116 28
rect 2892 -28 2948 -26
rect 4060 -26 4062 26
rect 4062 -26 4114 26
rect 4114 -26 4116 26
rect 5228 26 5284 28
rect 4060 -28 4116 -26
rect 5228 -26 5230 26
rect 5230 -26 5282 26
rect 5282 -26 5284 26
rect 6396 26 6452 28
rect 5228 -28 5284 -26
rect 6396 -26 6398 26
rect 6398 -26 6450 26
rect 6450 -26 6452 26
rect 7564 26 7620 28
rect 6396 -28 6452 -26
rect 7564 -26 7566 26
rect 7566 -26 7618 26
rect 7618 -26 7620 26
rect 8732 26 8788 28
rect 7564 -28 7620 -26
rect 8732 -26 8734 26
rect 8734 -26 8786 26
rect 8786 -26 8788 26
rect 8732 -28 8788 -26
<< metal3 >>
rect 535 1442 633 1463
rect 535 1386 556 1442
rect 612 1386 633 1442
rect 535 1365 633 1386
rect 1703 1442 1801 1463
rect 1703 1386 1724 1442
rect 1780 1386 1801 1442
rect 1703 1365 1801 1386
rect 2871 1442 2969 1463
rect 2871 1386 2892 1442
rect 2948 1386 2969 1442
rect 2871 1365 2969 1386
rect 4039 1442 4137 1463
rect 4039 1386 4060 1442
rect 4116 1386 4137 1442
rect 4039 1365 4137 1386
rect 5207 1442 5305 1463
rect 5207 1386 5228 1442
rect 5284 1386 5305 1442
rect 5207 1365 5305 1386
rect 6375 1442 6473 1463
rect 6375 1386 6396 1442
rect 6452 1386 6473 1442
rect 6375 1365 6473 1386
rect 7543 1442 7641 1463
rect 7543 1386 7564 1442
rect 7620 1386 7641 1442
rect 7543 1365 7641 1386
rect 8711 1442 8809 1463
rect 8711 1386 8732 1442
rect 8788 1386 8809 1442
rect 8711 1365 8809 1386
rect 363 338 429 341
rect 1531 338 1597 341
rect 2699 338 2765 341
rect 3867 338 3933 341
rect 5035 338 5101 341
rect 6203 338 6269 341
rect 7371 338 7437 341
rect 8539 338 8605 341
rect 0 336 9344 338
rect 0 280 368 336
rect 424 280 1536 336
rect 1592 280 2704 336
rect 2760 280 3872 336
rect 3928 280 5040 336
rect 5096 280 6208 336
rect 6264 280 7376 336
rect 7432 280 8544 336
rect 8600 280 9344 336
rect 0 278 9344 280
rect 363 275 429 278
rect 1531 275 1597 278
rect 2699 275 2765 278
rect 3867 275 3933 278
rect 5035 275 5101 278
rect 6203 275 6269 278
rect 7371 275 7437 278
rect 8539 275 8605 278
rect 535 28 633 49
rect 535 -28 556 28
rect 612 -28 633 28
rect 535 -49 633 -28
rect 1703 28 1801 49
rect 1703 -28 1724 28
rect 1780 -28 1801 28
rect 1703 -49 1801 -28
rect 2871 28 2969 49
rect 2871 -28 2892 28
rect 2948 -28 2969 28
rect 2871 -49 2969 -28
rect 4039 28 4137 49
rect 4039 -28 4060 28
rect 4116 -28 4137 28
rect 4039 -49 4137 -28
rect 5207 28 5305 49
rect 5207 -28 5228 28
rect 5284 -28 5305 28
rect 5207 -49 5305 -28
rect 6375 28 6473 49
rect 6375 -28 6396 28
rect 6452 -28 6473 28
rect 6375 -49 6473 -28
rect 7543 28 7641 49
rect 7543 -28 7564 28
rect 7620 -28 7641 28
rect 7543 -49 7641 -28
rect 8711 28 8809 49
rect 8711 -28 8732 28
rect 8788 -28 8809 28
rect 8711 -49 8809 -28
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 8539 0 1 271
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 7371 0 1 271
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 6203 0 1 271
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 5035 0 1 271
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 3867 0 1 271
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 2699 0 1 271
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 1531 0 1 271
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 363 0 1 271
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 8727 0 1 -37
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 8728 0 1 -32
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 8731 0 1 -33
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 8727 0 1 1377
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 8728 0 1 1382
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 8731 0 1 1381
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 7559 0 1 -37
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 7560 0 1 -32
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 7563 0 1 -33
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 7559 0 1 1377
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 7560 0 1 1382
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 7563 0 1 1381
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 6391 0 1 -37
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 6392 0 1 -32
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 6395 0 1 -33
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 6391 0 1 1377
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 6392 0 1 1382
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 6395 0 1 1381
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 5223 0 1 -37
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 5224 0 1 -32
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 5227 0 1 -33
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 5223 0 1 1377
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 5224 0 1 1382
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 5227 0 1 1381
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 4055 0 1 -37
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 4056 0 1 -32
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 4059 0 1 -33
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1634918361
transform 1 0 4055 0 1 1377
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 4056 0 1 1382
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 4059 0 1 1381
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1634918361
transform 1 0 2887 0 1 -37
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 2888 0 1 -32
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 2891 0 1 -33
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1634918361
transform 1 0 2887 0 1 1377
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 2888 0 1 1382
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 2891 0 1 1381
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1634918361
transform 1 0 1719 0 1 -37
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 1720 0 1 -32
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1634918361
transform 1 0 1723 0 1 -33
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1634918361
transform 1 0 1719 0 1 1377
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 1720 0 1 1382
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1634918361
transform 1 0 1723 0 1 1381
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1634918361
transform 1 0 551 0 1 -37
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 552 0 1 -32
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1634918361
transform 1 0 555 0 1 -33
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1634918361
transform 1 0 551 0 1 1377
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 552 0 1 1382
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1634918361
transform 1 0 555 0 1 1381
box 0 0 1 1
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1634918361
transform 1 0 8176 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_1
timestamp 1634918361
transform 1 0 7008 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_2
timestamp 1634918361
transform 1 0 5840 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_3
timestamp 1634918361
transform 1 0 4672 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_4
timestamp 1634918361
transform 1 0 3504 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_5
timestamp 1634918361
transform 1 0 2336 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_6
timestamp 1634918361
transform 1 0 1168 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_7
timestamp 1634918361
transform 1 0 0 0 1 0
box -36 -43 1204 1467
<< labels >>
rlabel metal3 s 8711 1365 8809 1463 4 vdd
port 1 nsew
rlabel metal3 s 4039 1365 4137 1463 4 vdd
port 1 nsew
rlabel metal3 s 6375 1365 6473 1463 4 vdd
port 1 nsew
rlabel metal3 s 1703 1365 1801 1463 4 vdd
port 1 nsew
rlabel metal3 s 7543 1365 7641 1463 4 vdd
port 1 nsew
rlabel metal3 s 535 1365 633 1463 4 vdd
port 1 nsew
rlabel metal3 s 2871 1365 2969 1463 4 vdd
port 1 nsew
rlabel metal3 s 5207 1365 5305 1463 4 vdd
port 1 nsew
rlabel metal3 s 8711 -49 8809 49 4 gnd
port 2 nsew
rlabel metal3 s 7543 -49 7641 49 4 gnd
port 2 nsew
rlabel metal3 s 1703 -49 1801 49 4 gnd
port 2 nsew
rlabel metal3 s 535 -49 633 49 4 gnd
port 2 nsew
rlabel metal3 s 6375 -49 6473 49 4 gnd
port 2 nsew
rlabel metal3 s 2871 -49 2969 49 4 gnd
port 2 nsew
rlabel metal3 s 5207 -49 5305 49 4 gnd
port 2 nsew
rlabel metal3 s 4039 -49 4137 49 4 gnd
port 2 nsew
rlabel metal2 s 137 538 203 590 4 din_0
port 3 nsew
rlabel metal2 s 1082 609 1148 661 4 dout_0
port 4 nsew
rlabel metal2 s 1305 538 1371 590 4 din_1
port 5 nsew
rlabel metal2 s 2250 609 2316 661 4 dout_1
port 6 nsew
rlabel metal2 s 2473 538 2539 590 4 din_2
port 7 nsew
rlabel metal2 s 3418 609 3484 661 4 dout_2
port 8 nsew
rlabel metal2 s 3641 538 3707 590 4 din_3
port 9 nsew
rlabel metal2 s 4586 609 4652 661 4 dout_3
port 10 nsew
rlabel metal2 s 4809 538 4875 590 4 din_4
port 11 nsew
rlabel metal2 s 5754 609 5820 661 4 dout_4
port 12 nsew
rlabel metal2 s 5977 538 6043 590 4 din_5
port 13 nsew
rlabel metal2 s 6922 609 6988 661 4 dout_5
port 14 nsew
rlabel metal2 s 7145 538 7211 590 4 din_6
port 15 nsew
rlabel metal2 s 8090 609 8156 661 4 dout_6
port 16 nsew
rlabel metal2 s 8313 538 8379 590 4 din_7
port 17 nsew
rlabel metal2 s 9258 609 9324 661 4 dout_7
port 18 nsew
rlabel metal3 s 0 278 9344 338 4 clk
port 19 nsew
<< properties >>
string FIXED_BBOX 8727 -37 8793 0
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1229134
string GDS_START 1217948
<< end >>
