magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1286 -1286 1436 1434
<< pwell >>
rect -26 -26 176 174
<< scnmos >>
rect 60 0 90 148
<< ndiff >>
rect 0 91 60 148
rect 0 57 8 91
rect 42 57 60 91
rect 0 0 60 57
rect 90 0 150 148
<< ndiffc >>
rect 8 57 42 91
<< poly >>
rect 60 148 90 174
rect 60 -26 90 0
<< locali >>
rect 8 91 42 107
rect 8 41 42 57
use contact_11  contact_11_0
timestamp 1634918361
transform 1 0 0 0 1 41
box 0 0 1 1
<< labels >>
rlabel poly s 75 74 75 74 4 G
port 1 nsew
rlabel locali s 25 74 25 74 4 S
port 2 nsew
rlabel mvpsubdiff s 125 74 125 74 4 D
<< properties >>
string FIXED_BBOX -25 -26 175 174
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 879296
string GDS_START 878608
<< end >>
