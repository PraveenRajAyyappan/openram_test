magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 806130
string GDS_START 805806
<< end >>
