magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1296 -1277 2690 2731
<< locali >>
rect 0 1397 1394 1431
rect 330 708 364 1151
rect 330 674 459 708
rect 883 674 917 708
rect 212 485 246 551
rect 112 237 146 303
rect 0 -17 1394 17
use pdriver_0  pdriver_0_0
timestamp 1634918361
transform 1 0 378 0 1 0
box -36 -17 1052 1471
use pnand2_0  pnand2_0_0
timestamp 1634918361
transform 1 0 0 0 1 0
box -36 -17 414 1471
<< labels >>
rlabel locali s 900 691 900 691 4 Z
port 1 nsew
rlabel locali s 129 270 129 270 4 A
port 2 nsew
rlabel locali s 229 518 229 518 4 B
port 3 nsew
rlabel locali s 697 0 697 0 4 gnd
port 4 nsew
rlabel locali s 697 1414 697 1414 4 vdd
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1394 1414
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1112076
string GDS_START 1111002
<< end >>
