magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1296 -1277 3006 2731
<< locali >>
rect 0 1397 1710 1431
rect 430 724 464 1167
rect 430 690 559 724
rect 1091 690 1125 724
rect 345 485 379 551
rect 212 361 246 427
rect 79 237 113 303
rect 0 -17 1710 17
use pdriver_3  pdriver_3_0
timestamp 1634918361
transform 1 0 478 0 1 0
box -36 -17 1268 1471
use pnand3  pnand3_0
timestamp 1634918361
transform 1 0 0 0 1 0
box -36 -17 514 1471
<< labels >>
rlabel locali s 1108 707 1108 707 4 Z
port 1 nsew
rlabel locali s 96 270 96 270 4 A
port 2 nsew
rlabel locali s 229 394 229 394 4 B
port 3 nsew
rlabel locali s 362 518 362 518 4 C
port 4 nsew
rlabel locali s 855 0 855 0 4 gnd
port 5 nsew
rlabel locali s 855 1414 855 1414 4 vdd
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 1710 1414
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1128118
string GDS_START 1126938
<< end >>
