magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1335 -1309 3136 14043
<< locali >>
rect 639 12743 673 12759
rect 639 12693 673 12709
rect 1375 12743 1409 12759
rect 1375 12693 1409 12709
rect 64 11998 98 12014
rect 64 11948 98 11964
rect 179 11998 213 12014
rect 179 11948 213 11964
rect 432 11998 466 12014
rect 432 11948 466 11964
rect 800 11998 834 12014
rect 800 11948 834 11964
rect 1168 11998 1202 12014
rect 1168 11948 1202 11964
rect 1536 11998 1570 12014
rect 1536 11948 1570 11964
rect 639 11329 673 11345
rect 639 11279 673 11295
rect 1375 11329 1409 11345
rect 1375 11279 1409 11295
rect 64 10660 98 10676
rect 64 10610 98 10626
rect 179 10660 213 10676
rect 179 10610 213 10626
rect 432 10660 466 10676
rect 432 10610 466 10626
rect 800 10660 834 10676
rect 800 10610 834 10626
rect 1168 10660 1202 10676
rect 1168 10610 1202 10626
rect 1536 10660 1570 10676
rect 1536 10610 1570 10626
rect 639 9915 673 9931
rect 639 9865 673 9881
rect 1375 9915 1409 9931
rect 1375 9865 1409 9881
rect 64 9170 98 9186
rect 64 9120 98 9136
rect 179 9170 213 9186
rect 179 9120 213 9136
rect 432 9170 466 9186
rect 432 9120 466 9136
rect 800 9170 834 9186
rect 800 9120 834 9136
rect 1168 9170 1202 9186
rect 1168 9120 1202 9136
rect 1536 9170 1570 9186
rect 1536 9120 1570 9136
rect 639 8501 673 8517
rect 639 8451 673 8467
rect 1375 8501 1409 8517
rect 1375 8451 1409 8467
rect 64 7832 98 7848
rect 64 7782 98 7798
rect 179 7832 213 7848
rect 179 7782 213 7798
rect 432 7832 466 7848
rect 432 7782 466 7798
rect 800 7832 834 7848
rect 800 7782 834 7798
rect 1168 7832 1202 7848
rect 1168 7782 1202 7798
rect 1536 7832 1570 7848
rect 1536 7782 1570 7798
rect 639 7087 673 7103
rect 639 7037 673 7053
rect 1375 7087 1409 7103
rect 1375 7037 1409 7053
rect 64 6342 98 6358
rect 64 6292 98 6308
rect 179 6342 213 6358
rect 179 6292 213 6308
rect 432 6342 466 6358
rect 432 6292 466 6308
rect 800 6342 834 6358
rect 800 6292 834 6308
rect 1168 6342 1202 6358
rect 1168 6292 1202 6308
rect 1536 6342 1570 6358
rect 1536 6292 1570 6308
rect 639 5673 673 5689
rect 639 5623 673 5639
rect 1375 5673 1409 5689
rect 1375 5623 1409 5639
rect 64 5004 98 5020
rect 64 4954 98 4970
rect 179 5004 213 5020
rect 179 4954 213 4970
rect 432 5004 466 5020
rect 432 4954 466 4970
rect 800 5004 834 5020
rect 800 4954 834 4970
rect 1168 5004 1202 5020
rect 1168 4954 1202 4970
rect 1536 5004 1570 5020
rect 1536 4954 1570 4970
rect 639 4259 673 4275
rect 639 4209 673 4225
rect 1375 4259 1409 4275
rect 1375 4209 1409 4225
rect 64 3514 98 3530
rect 64 3464 98 3480
rect 179 3514 213 3530
rect 179 3464 213 3480
rect 432 3514 466 3530
rect 432 3464 466 3480
rect 800 3514 834 3530
rect 800 3464 834 3480
rect 1168 3514 1202 3530
rect 1168 3464 1202 3480
rect 1536 3514 1570 3530
rect 1536 3464 1570 3480
rect 639 2845 673 2861
rect 639 2795 673 2811
rect 1375 2845 1409 2861
rect 1375 2795 1409 2811
rect 64 2176 98 2192
rect 64 2126 98 2142
rect 179 2176 213 2192
rect 179 2126 213 2142
rect 432 2176 466 2192
rect 432 2126 466 2142
rect 800 2176 834 2192
rect 800 2126 834 2142
rect 1168 2176 1202 2192
rect 1168 2126 1202 2142
rect 1536 2176 1570 2192
rect 1536 2126 1570 2142
rect 639 1431 673 1447
rect 639 1381 673 1397
rect 1375 1431 1409 1447
rect 1375 1381 1409 1397
rect -60 686 -26 702
rect 64 686 98 702
rect -26 652 64 686
rect -60 636 -26 652
rect 64 636 98 652
rect 179 686 213 702
rect 179 636 213 652
rect 432 686 466 702
rect 432 636 466 652
rect 800 686 834 702
rect 800 636 834 652
rect 1168 686 1202 702
rect 1168 636 1202 652
rect 1536 686 1570 702
rect 1536 636 1570 652
rect 639 17 673 33
rect 639 -33 673 -17
rect 1375 17 1409 33
rect 1375 -33 1409 -17
<< viali >>
rect 639 12709 673 12743
rect 1375 12709 1409 12743
rect 64 11964 98 11998
rect 179 11964 213 11998
rect 432 11964 466 11998
rect 800 11964 834 11998
rect 1168 11964 1202 11998
rect 1536 11964 1570 11998
rect 639 11295 673 11329
rect 1375 11295 1409 11329
rect 64 10626 98 10660
rect 179 10626 213 10660
rect 432 10626 466 10660
rect 800 10626 834 10660
rect 1168 10626 1202 10660
rect 1536 10626 1570 10660
rect 639 9881 673 9915
rect 1375 9881 1409 9915
rect 64 9136 98 9170
rect 179 9136 213 9170
rect 432 9136 466 9170
rect 800 9136 834 9170
rect 1168 9136 1202 9170
rect 1536 9136 1570 9170
rect 639 8467 673 8501
rect 1375 8467 1409 8501
rect 64 7798 98 7832
rect 179 7798 213 7832
rect 432 7798 466 7832
rect 800 7798 834 7832
rect 1168 7798 1202 7832
rect 1536 7798 1570 7832
rect 639 7053 673 7087
rect 1375 7053 1409 7087
rect 64 6308 98 6342
rect 179 6308 213 6342
rect 432 6308 466 6342
rect 800 6308 834 6342
rect 1168 6308 1202 6342
rect 1536 6308 1570 6342
rect 639 5639 673 5673
rect 1375 5639 1409 5673
rect 64 4970 98 5004
rect 179 4970 213 5004
rect 432 4970 466 5004
rect 800 4970 834 5004
rect 1168 4970 1202 5004
rect 1536 4970 1570 5004
rect 639 4225 673 4259
rect 1375 4225 1409 4259
rect 64 3480 98 3514
rect 179 3480 213 3514
rect 432 3480 466 3514
rect 800 3480 834 3514
rect 1168 3480 1202 3514
rect 1536 3480 1570 3514
rect 639 2811 673 2845
rect 1375 2811 1409 2845
rect 64 2142 98 2176
rect 179 2142 213 2176
rect 432 2142 466 2176
rect 800 2142 834 2176
rect 1168 2142 1202 2176
rect 1536 2142 1570 2176
rect 639 1397 673 1431
rect 1375 1397 1409 1431
rect -60 652 -26 686
rect 64 652 98 686
rect 179 652 213 686
rect 432 652 466 686
rect 800 652 834 686
rect 1168 652 1202 686
rect 1536 652 1570 686
rect 639 -17 673 17
rect 1375 -17 1409 17
<< metal1 >>
rect 624 12700 630 12752
rect 682 12700 688 12752
rect 1360 12700 1366 12752
rect 1418 12700 1424 12752
rect 49 11955 55 12007
rect 107 11955 113 12007
rect 164 11955 170 12007
rect 222 11955 228 12007
rect 417 11955 423 12007
rect 475 11955 481 12007
rect 785 11955 791 12007
rect 843 11955 849 12007
rect 1153 11955 1159 12007
rect 1211 11955 1217 12007
rect 1521 11955 1527 12007
rect 1579 11955 1585 12007
rect 624 11286 630 11338
rect 682 11286 688 11338
rect 1360 11286 1366 11338
rect 1418 11286 1424 11338
rect 49 10617 55 10669
rect 107 10617 113 10669
rect 164 10617 170 10669
rect 222 10617 228 10669
rect 417 10617 423 10669
rect 475 10617 481 10669
rect 785 10617 791 10669
rect 843 10617 849 10669
rect 1153 10617 1159 10669
rect 1211 10617 1217 10669
rect 1521 10617 1527 10669
rect 1579 10617 1585 10669
rect 624 9872 630 9924
rect 682 9872 688 9924
rect 1360 9872 1366 9924
rect 1418 9872 1424 9924
rect 49 9127 55 9179
rect 107 9127 113 9179
rect 164 9127 170 9179
rect 222 9127 228 9179
rect 417 9127 423 9179
rect 475 9127 481 9179
rect 785 9127 791 9179
rect 843 9127 849 9179
rect 1153 9127 1159 9179
rect 1211 9127 1217 9179
rect 1521 9127 1527 9179
rect 1579 9127 1585 9179
rect 624 8458 630 8510
rect 682 8458 688 8510
rect 1360 8458 1366 8510
rect 1418 8458 1424 8510
rect 49 7789 55 7841
rect 107 7789 113 7841
rect 164 7789 170 7841
rect 222 7789 228 7841
rect 417 7789 423 7841
rect 475 7789 481 7841
rect 785 7789 791 7841
rect 843 7789 849 7841
rect 1153 7789 1159 7841
rect 1211 7789 1217 7841
rect 1521 7789 1527 7841
rect 1579 7789 1585 7841
rect 624 7044 630 7096
rect 682 7044 688 7096
rect 1360 7044 1366 7096
rect 1418 7044 1424 7096
rect 49 6299 55 6351
rect 107 6299 113 6351
rect 164 6299 170 6351
rect 222 6299 228 6351
rect 417 6299 423 6351
rect 475 6299 481 6351
rect 785 6299 791 6351
rect 843 6299 849 6351
rect 1153 6299 1159 6351
rect 1211 6299 1217 6351
rect 1521 6299 1527 6351
rect 1579 6299 1585 6351
rect 624 5630 630 5682
rect 682 5630 688 5682
rect 1360 5630 1366 5682
rect 1418 5630 1424 5682
rect 49 4961 55 5013
rect 107 4961 113 5013
rect 164 4961 170 5013
rect 222 4961 228 5013
rect 417 4961 423 5013
rect 475 4961 481 5013
rect 785 4961 791 5013
rect 843 4961 849 5013
rect 1153 4961 1159 5013
rect 1211 4961 1217 5013
rect 1521 4961 1527 5013
rect 1579 4961 1585 5013
rect 624 4216 630 4268
rect 682 4216 688 4268
rect 1360 4216 1366 4268
rect 1418 4216 1424 4268
rect 49 3471 55 3523
rect 107 3471 113 3523
rect 164 3471 170 3523
rect 222 3471 228 3523
rect 417 3471 423 3523
rect 475 3471 481 3523
rect 785 3471 791 3523
rect 843 3471 849 3523
rect 1153 3471 1159 3523
rect 1211 3471 1217 3523
rect 1521 3471 1527 3523
rect 1579 3471 1585 3523
rect 624 2802 630 2854
rect 682 2802 688 2854
rect 1360 2802 1366 2854
rect 1418 2802 1424 2854
rect 49 2133 55 2185
rect 107 2133 113 2185
rect 164 2133 170 2185
rect 222 2133 228 2185
rect 417 2133 423 2185
rect 475 2133 481 2185
rect 785 2133 791 2185
rect 843 2133 849 2185
rect 1153 2133 1159 2185
rect 1211 2133 1217 2185
rect 1521 2133 1527 2185
rect 1579 2133 1585 2185
rect 624 1388 630 1440
rect 682 1388 688 1440
rect 1360 1388 1366 1440
rect 1418 1388 1424 1440
rect -75 643 -69 695
rect -17 643 -11 695
rect 49 643 55 695
rect 107 643 113 695
rect 164 643 170 695
rect 222 643 228 695
rect 417 643 423 695
rect 475 643 481 695
rect 785 643 791 695
rect 843 643 849 695
rect 1153 643 1159 695
rect 1211 643 1217 695
rect 1521 643 1527 695
rect 1579 643 1585 695
rect 624 -26 630 26
rect 682 -26 688 26
rect 1360 -26 1366 26
rect 1418 -26 1424 26
<< via1 >>
rect 630 12743 682 12752
rect 630 12709 639 12743
rect 639 12709 673 12743
rect 673 12709 682 12743
rect 630 12700 682 12709
rect 1366 12743 1418 12752
rect 1366 12709 1375 12743
rect 1375 12709 1409 12743
rect 1409 12709 1418 12743
rect 1366 12700 1418 12709
rect 55 11998 107 12007
rect 55 11964 64 11998
rect 64 11964 98 11998
rect 98 11964 107 11998
rect 55 11955 107 11964
rect 170 11998 222 12007
rect 170 11964 179 11998
rect 179 11964 213 11998
rect 213 11964 222 11998
rect 170 11955 222 11964
rect 423 11998 475 12007
rect 423 11964 432 11998
rect 432 11964 466 11998
rect 466 11964 475 11998
rect 423 11955 475 11964
rect 791 11998 843 12007
rect 791 11964 800 11998
rect 800 11964 834 11998
rect 834 11964 843 11998
rect 791 11955 843 11964
rect 1159 11998 1211 12007
rect 1159 11964 1168 11998
rect 1168 11964 1202 11998
rect 1202 11964 1211 11998
rect 1159 11955 1211 11964
rect 1527 11998 1579 12007
rect 1527 11964 1536 11998
rect 1536 11964 1570 11998
rect 1570 11964 1579 11998
rect 1527 11955 1579 11964
rect 630 11329 682 11338
rect 630 11295 639 11329
rect 639 11295 673 11329
rect 673 11295 682 11329
rect 630 11286 682 11295
rect 1366 11329 1418 11338
rect 1366 11295 1375 11329
rect 1375 11295 1409 11329
rect 1409 11295 1418 11329
rect 1366 11286 1418 11295
rect 55 10660 107 10669
rect 55 10626 64 10660
rect 64 10626 98 10660
rect 98 10626 107 10660
rect 55 10617 107 10626
rect 170 10660 222 10669
rect 170 10626 179 10660
rect 179 10626 213 10660
rect 213 10626 222 10660
rect 170 10617 222 10626
rect 423 10660 475 10669
rect 423 10626 432 10660
rect 432 10626 466 10660
rect 466 10626 475 10660
rect 423 10617 475 10626
rect 791 10660 843 10669
rect 791 10626 800 10660
rect 800 10626 834 10660
rect 834 10626 843 10660
rect 791 10617 843 10626
rect 1159 10660 1211 10669
rect 1159 10626 1168 10660
rect 1168 10626 1202 10660
rect 1202 10626 1211 10660
rect 1159 10617 1211 10626
rect 1527 10660 1579 10669
rect 1527 10626 1536 10660
rect 1536 10626 1570 10660
rect 1570 10626 1579 10660
rect 1527 10617 1579 10626
rect 630 9915 682 9924
rect 630 9881 639 9915
rect 639 9881 673 9915
rect 673 9881 682 9915
rect 630 9872 682 9881
rect 1366 9915 1418 9924
rect 1366 9881 1375 9915
rect 1375 9881 1409 9915
rect 1409 9881 1418 9915
rect 1366 9872 1418 9881
rect 55 9170 107 9179
rect 55 9136 64 9170
rect 64 9136 98 9170
rect 98 9136 107 9170
rect 55 9127 107 9136
rect 170 9170 222 9179
rect 170 9136 179 9170
rect 179 9136 213 9170
rect 213 9136 222 9170
rect 170 9127 222 9136
rect 423 9170 475 9179
rect 423 9136 432 9170
rect 432 9136 466 9170
rect 466 9136 475 9170
rect 423 9127 475 9136
rect 791 9170 843 9179
rect 791 9136 800 9170
rect 800 9136 834 9170
rect 834 9136 843 9170
rect 791 9127 843 9136
rect 1159 9170 1211 9179
rect 1159 9136 1168 9170
rect 1168 9136 1202 9170
rect 1202 9136 1211 9170
rect 1159 9127 1211 9136
rect 1527 9170 1579 9179
rect 1527 9136 1536 9170
rect 1536 9136 1570 9170
rect 1570 9136 1579 9170
rect 1527 9127 1579 9136
rect 630 8501 682 8510
rect 630 8467 639 8501
rect 639 8467 673 8501
rect 673 8467 682 8501
rect 630 8458 682 8467
rect 1366 8501 1418 8510
rect 1366 8467 1375 8501
rect 1375 8467 1409 8501
rect 1409 8467 1418 8501
rect 1366 8458 1418 8467
rect 55 7832 107 7841
rect 55 7798 64 7832
rect 64 7798 98 7832
rect 98 7798 107 7832
rect 55 7789 107 7798
rect 170 7832 222 7841
rect 170 7798 179 7832
rect 179 7798 213 7832
rect 213 7798 222 7832
rect 170 7789 222 7798
rect 423 7832 475 7841
rect 423 7798 432 7832
rect 432 7798 466 7832
rect 466 7798 475 7832
rect 423 7789 475 7798
rect 791 7832 843 7841
rect 791 7798 800 7832
rect 800 7798 834 7832
rect 834 7798 843 7832
rect 791 7789 843 7798
rect 1159 7832 1211 7841
rect 1159 7798 1168 7832
rect 1168 7798 1202 7832
rect 1202 7798 1211 7832
rect 1159 7789 1211 7798
rect 1527 7832 1579 7841
rect 1527 7798 1536 7832
rect 1536 7798 1570 7832
rect 1570 7798 1579 7832
rect 1527 7789 1579 7798
rect 630 7087 682 7096
rect 630 7053 639 7087
rect 639 7053 673 7087
rect 673 7053 682 7087
rect 630 7044 682 7053
rect 1366 7087 1418 7096
rect 1366 7053 1375 7087
rect 1375 7053 1409 7087
rect 1409 7053 1418 7087
rect 1366 7044 1418 7053
rect 55 6342 107 6351
rect 55 6308 64 6342
rect 64 6308 98 6342
rect 98 6308 107 6342
rect 55 6299 107 6308
rect 170 6342 222 6351
rect 170 6308 179 6342
rect 179 6308 213 6342
rect 213 6308 222 6342
rect 170 6299 222 6308
rect 423 6342 475 6351
rect 423 6308 432 6342
rect 432 6308 466 6342
rect 466 6308 475 6342
rect 423 6299 475 6308
rect 791 6342 843 6351
rect 791 6308 800 6342
rect 800 6308 834 6342
rect 834 6308 843 6342
rect 791 6299 843 6308
rect 1159 6342 1211 6351
rect 1159 6308 1168 6342
rect 1168 6308 1202 6342
rect 1202 6308 1211 6342
rect 1159 6299 1211 6308
rect 1527 6342 1579 6351
rect 1527 6308 1536 6342
rect 1536 6308 1570 6342
rect 1570 6308 1579 6342
rect 1527 6299 1579 6308
rect 630 5673 682 5682
rect 630 5639 639 5673
rect 639 5639 673 5673
rect 673 5639 682 5673
rect 630 5630 682 5639
rect 1366 5673 1418 5682
rect 1366 5639 1375 5673
rect 1375 5639 1409 5673
rect 1409 5639 1418 5673
rect 1366 5630 1418 5639
rect 55 5004 107 5013
rect 55 4970 64 5004
rect 64 4970 98 5004
rect 98 4970 107 5004
rect 55 4961 107 4970
rect 170 5004 222 5013
rect 170 4970 179 5004
rect 179 4970 213 5004
rect 213 4970 222 5004
rect 170 4961 222 4970
rect 423 5004 475 5013
rect 423 4970 432 5004
rect 432 4970 466 5004
rect 466 4970 475 5004
rect 423 4961 475 4970
rect 791 5004 843 5013
rect 791 4970 800 5004
rect 800 4970 834 5004
rect 834 4970 843 5004
rect 791 4961 843 4970
rect 1159 5004 1211 5013
rect 1159 4970 1168 5004
rect 1168 4970 1202 5004
rect 1202 4970 1211 5004
rect 1159 4961 1211 4970
rect 1527 5004 1579 5013
rect 1527 4970 1536 5004
rect 1536 4970 1570 5004
rect 1570 4970 1579 5004
rect 1527 4961 1579 4970
rect 630 4259 682 4268
rect 630 4225 639 4259
rect 639 4225 673 4259
rect 673 4225 682 4259
rect 630 4216 682 4225
rect 1366 4259 1418 4268
rect 1366 4225 1375 4259
rect 1375 4225 1409 4259
rect 1409 4225 1418 4259
rect 1366 4216 1418 4225
rect 55 3514 107 3523
rect 55 3480 64 3514
rect 64 3480 98 3514
rect 98 3480 107 3514
rect 55 3471 107 3480
rect 170 3514 222 3523
rect 170 3480 179 3514
rect 179 3480 213 3514
rect 213 3480 222 3514
rect 170 3471 222 3480
rect 423 3514 475 3523
rect 423 3480 432 3514
rect 432 3480 466 3514
rect 466 3480 475 3514
rect 423 3471 475 3480
rect 791 3514 843 3523
rect 791 3480 800 3514
rect 800 3480 834 3514
rect 834 3480 843 3514
rect 791 3471 843 3480
rect 1159 3514 1211 3523
rect 1159 3480 1168 3514
rect 1168 3480 1202 3514
rect 1202 3480 1211 3514
rect 1159 3471 1211 3480
rect 1527 3514 1579 3523
rect 1527 3480 1536 3514
rect 1536 3480 1570 3514
rect 1570 3480 1579 3514
rect 1527 3471 1579 3480
rect 630 2845 682 2854
rect 630 2811 639 2845
rect 639 2811 673 2845
rect 673 2811 682 2845
rect 630 2802 682 2811
rect 1366 2845 1418 2854
rect 1366 2811 1375 2845
rect 1375 2811 1409 2845
rect 1409 2811 1418 2845
rect 1366 2802 1418 2811
rect 55 2176 107 2185
rect 55 2142 64 2176
rect 64 2142 98 2176
rect 98 2142 107 2176
rect 55 2133 107 2142
rect 170 2176 222 2185
rect 170 2142 179 2176
rect 179 2142 213 2176
rect 213 2142 222 2176
rect 170 2133 222 2142
rect 423 2176 475 2185
rect 423 2142 432 2176
rect 432 2142 466 2176
rect 466 2142 475 2176
rect 423 2133 475 2142
rect 791 2176 843 2185
rect 791 2142 800 2176
rect 800 2142 834 2176
rect 834 2142 843 2176
rect 791 2133 843 2142
rect 1159 2176 1211 2185
rect 1159 2142 1168 2176
rect 1168 2142 1202 2176
rect 1202 2142 1211 2176
rect 1159 2133 1211 2142
rect 1527 2176 1579 2185
rect 1527 2142 1536 2176
rect 1536 2142 1570 2176
rect 1570 2142 1579 2176
rect 1527 2133 1579 2142
rect 630 1431 682 1440
rect 630 1397 639 1431
rect 639 1397 673 1431
rect 673 1397 682 1431
rect 630 1388 682 1397
rect 1366 1431 1418 1440
rect 1366 1397 1375 1431
rect 1375 1397 1409 1431
rect 1409 1397 1418 1431
rect 1366 1388 1418 1397
rect -69 686 -17 695
rect -69 652 -60 686
rect -60 652 -26 686
rect -26 652 -17 686
rect -69 643 -17 652
rect 55 686 107 695
rect 55 652 64 686
rect 64 652 98 686
rect 98 652 107 686
rect 55 643 107 652
rect 170 686 222 695
rect 170 652 179 686
rect 179 652 213 686
rect 213 652 222 686
rect 170 643 222 652
rect 423 686 475 695
rect 423 652 432 686
rect 432 652 466 686
rect 466 652 475 686
rect 423 643 475 652
rect 791 686 843 695
rect 791 652 800 686
rect 800 652 834 686
rect 834 652 843 686
rect 791 643 843 652
rect 1159 686 1211 695
rect 1159 652 1168 686
rect 1168 652 1202 686
rect 1202 652 1211 686
rect 1159 643 1211 652
rect 1527 686 1579 695
rect 1527 652 1536 686
rect 1536 652 1570 686
rect 1570 652 1579 686
rect 1527 643 1579 652
rect 630 17 682 26
rect 630 -17 639 17
rect 639 -17 673 17
rect 673 -17 682 17
rect 630 -26 682 -17
rect 1366 17 1418 26
rect 1366 -17 1375 17
rect 1375 -17 1409 17
rect 1409 -17 1418 17
rect 1366 -26 1418 -17
<< metal2 >>
rect 628 12754 684 12763
rect 628 12689 684 12698
rect 1364 12754 1420 12763
rect 1364 12689 1420 12698
rect 55 12007 107 12013
rect 55 11949 107 11955
rect 168 12009 224 12018
rect 67 11326 95 11949
rect 168 11944 224 11953
rect 421 12009 477 12018
rect 421 11944 477 11953
rect 789 12009 845 12018
rect 789 11944 845 11953
rect 1157 12009 1213 12018
rect 1157 11944 1213 11953
rect 1525 12009 1581 12018
rect 1525 11944 1581 11953
rect 628 11340 684 11349
rect 67 11298 210 11326
rect 182 10680 210 11298
rect 628 11275 684 11284
rect 1364 11340 1420 11349
rect 1364 11275 1420 11284
rect 55 10669 107 10675
rect 55 10611 107 10617
rect 168 10671 224 10680
rect 67 9912 95 10611
rect 168 10606 224 10615
rect 421 10671 477 10680
rect 421 10606 477 10615
rect 789 10671 845 10680
rect 789 10606 845 10615
rect 1157 10671 1213 10680
rect 1157 10606 1213 10615
rect 1525 10671 1581 10680
rect 1525 10606 1581 10615
rect 628 9926 684 9935
rect 67 9884 210 9912
rect 182 9190 210 9884
rect 628 9861 684 9870
rect 1364 9926 1420 9935
rect 1364 9861 1420 9870
rect 55 9179 107 9185
rect 55 9121 107 9127
rect 168 9181 224 9190
rect 67 8498 95 9121
rect 168 9116 224 9125
rect 421 9181 477 9190
rect 421 9116 477 9125
rect 789 9181 845 9190
rect 789 9116 845 9125
rect 1157 9181 1213 9190
rect 1157 9116 1213 9125
rect 1525 9181 1581 9190
rect 1525 9116 1581 9125
rect 628 8512 684 8521
rect 67 8470 210 8498
rect 182 7852 210 8470
rect 628 8447 684 8456
rect 1364 8512 1420 8521
rect 1364 8447 1420 8456
rect 55 7841 107 7847
rect 55 7783 107 7789
rect 168 7843 224 7852
rect 67 7084 95 7783
rect 168 7778 224 7787
rect 421 7843 477 7852
rect 421 7778 477 7787
rect 789 7843 845 7852
rect 789 7778 845 7787
rect 1157 7843 1213 7852
rect 1157 7778 1213 7787
rect 1525 7843 1581 7852
rect 1525 7778 1581 7787
rect 628 7098 684 7107
rect 67 7056 210 7084
rect 182 6362 210 7056
rect 628 7033 684 7042
rect 1364 7098 1420 7107
rect 1364 7033 1420 7042
rect 55 6351 107 6357
rect 55 6293 107 6299
rect 168 6353 224 6362
rect 67 5670 95 6293
rect 168 6288 224 6297
rect 421 6353 477 6362
rect 421 6288 477 6297
rect 789 6353 845 6362
rect 789 6288 845 6297
rect 1157 6353 1213 6362
rect 1157 6288 1213 6297
rect 1525 6353 1581 6362
rect 1525 6288 1581 6297
rect 628 5684 684 5693
rect 67 5642 210 5670
rect 182 5024 210 5642
rect 628 5619 684 5628
rect 1364 5684 1420 5693
rect 1364 5619 1420 5628
rect 55 5013 107 5019
rect 55 4955 107 4961
rect 168 5015 224 5024
rect 67 4256 95 4955
rect 168 4950 224 4959
rect 421 5015 477 5024
rect 421 4950 477 4959
rect 789 5015 845 5024
rect 789 4950 845 4959
rect 1157 5015 1213 5024
rect 1157 4950 1213 4959
rect 1525 5015 1581 5024
rect 1525 4950 1581 4959
rect 628 4270 684 4279
rect 67 4228 210 4256
rect 182 3534 210 4228
rect 628 4205 684 4214
rect 1364 4270 1420 4279
rect 1364 4205 1420 4214
rect 55 3523 107 3529
rect 55 3465 107 3471
rect 168 3525 224 3534
rect 67 2842 95 3465
rect 168 3460 224 3469
rect 421 3525 477 3534
rect 421 3460 477 3469
rect 789 3525 845 3534
rect 789 3460 845 3469
rect 1157 3525 1213 3534
rect 1157 3460 1213 3469
rect 1525 3525 1581 3534
rect 1525 3460 1581 3469
rect 628 2856 684 2865
rect 67 2814 210 2842
rect 182 2196 210 2814
rect 628 2791 684 2800
rect 1364 2856 1420 2865
rect 1364 2791 1420 2800
rect 55 2185 107 2191
rect 55 2127 107 2133
rect 168 2187 224 2196
rect 67 1428 95 2127
rect 168 2122 224 2131
rect 421 2187 477 2196
rect 421 2122 477 2131
rect 789 2187 845 2196
rect 789 2122 845 2131
rect 1157 2187 1213 2196
rect 1157 2122 1213 2131
rect 1525 2187 1581 2196
rect 1525 2122 1581 2131
rect 628 1442 684 1451
rect 67 1400 210 1428
rect 182 706 210 1400
rect 628 1377 684 1386
rect 1364 1442 1420 1451
rect 1364 1377 1420 1386
rect -69 695 -17 701
rect -69 637 -17 643
rect 55 695 107 701
rect 55 637 107 643
rect 168 697 224 706
rect 168 632 224 641
rect 421 697 477 706
rect 421 632 477 641
rect 789 697 845 706
rect 789 632 845 641
rect 1157 697 1213 706
rect 1157 632 1213 641
rect 1525 697 1581 706
rect 1525 632 1581 641
rect 628 28 684 37
rect 628 -37 684 -28
rect 1364 28 1420 37
rect 1364 -37 1420 -28
<< via2 >>
rect 628 12752 684 12754
rect 628 12700 630 12752
rect 630 12700 682 12752
rect 682 12700 684 12752
rect 628 12698 684 12700
rect 1364 12752 1420 12754
rect 1364 12700 1366 12752
rect 1366 12700 1418 12752
rect 1418 12700 1420 12752
rect 1364 12698 1420 12700
rect 168 12007 224 12009
rect 168 11955 170 12007
rect 170 11955 222 12007
rect 222 11955 224 12007
rect 168 11953 224 11955
rect 421 12007 477 12009
rect 421 11955 423 12007
rect 423 11955 475 12007
rect 475 11955 477 12007
rect 421 11953 477 11955
rect 789 12007 845 12009
rect 789 11955 791 12007
rect 791 11955 843 12007
rect 843 11955 845 12007
rect 789 11953 845 11955
rect 1157 12007 1213 12009
rect 1157 11955 1159 12007
rect 1159 11955 1211 12007
rect 1211 11955 1213 12007
rect 1157 11953 1213 11955
rect 1525 12007 1581 12009
rect 1525 11955 1527 12007
rect 1527 11955 1579 12007
rect 1579 11955 1581 12007
rect 1525 11953 1581 11955
rect 628 11338 684 11340
rect 628 11286 630 11338
rect 630 11286 682 11338
rect 682 11286 684 11338
rect 628 11284 684 11286
rect 1364 11338 1420 11340
rect 1364 11286 1366 11338
rect 1366 11286 1418 11338
rect 1418 11286 1420 11338
rect 1364 11284 1420 11286
rect 168 10669 224 10671
rect 168 10617 170 10669
rect 170 10617 222 10669
rect 222 10617 224 10669
rect 168 10615 224 10617
rect 421 10669 477 10671
rect 421 10617 423 10669
rect 423 10617 475 10669
rect 475 10617 477 10669
rect 421 10615 477 10617
rect 789 10669 845 10671
rect 789 10617 791 10669
rect 791 10617 843 10669
rect 843 10617 845 10669
rect 789 10615 845 10617
rect 1157 10669 1213 10671
rect 1157 10617 1159 10669
rect 1159 10617 1211 10669
rect 1211 10617 1213 10669
rect 1157 10615 1213 10617
rect 1525 10669 1581 10671
rect 1525 10617 1527 10669
rect 1527 10617 1579 10669
rect 1579 10617 1581 10669
rect 1525 10615 1581 10617
rect 628 9924 684 9926
rect 628 9872 630 9924
rect 630 9872 682 9924
rect 682 9872 684 9924
rect 628 9870 684 9872
rect 1364 9924 1420 9926
rect 1364 9872 1366 9924
rect 1366 9872 1418 9924
rect 1418 9872 1420 9924
rect 1364 9870 1420 9872
rect 168 9179 224 9181
rect 168 9127 170 9179
rect 170 9127 222 9179
rect 222 9127 224 9179
rect 168 9125 224 9127
rect 421 9179 477 9181
rect 421 9127 423 9179
rect 423 9127 475 9179
rect 475 9127 477 9179
rect 421 9125 477 9127
rect 789 9179 845 9181
rect 789 9127 791 9179
rect 791 9127 843 9179
rect 843 9127 845 9179
rect 789 9125 845 9127
rect 1157 9179 1213 9181
rect 1157 9127 1159 9179
rect 1159 9127 1211 9179
rect 1211 9127 1213 9179
rect 1157 9125 1213 9127
rect 1525 9179 1581 9181
rect 1525 9127 1527 9179
rect 1527 9127 1579 9179
rect 1579 9127 1581 9179
rect 1525 9125 1581 9127
rect 628 8510 684 8512
rect 628 8458 630 8510
rect 630 8458 682 8510
rect 682 8458 684 8510
rect 628 8456 684 8458
rect 1364 8510 1420 8512
rect 1364 8458 1366 8510
rect 1366 8458 1418 8510
rect 1418 8458 1420 8510
rect 1364 8456 1420 8458
rect 168 7841 224 7843
rect 168 7789 170 7841
rect 170 7789 222 7841
rect 222 7789 224 7841
rect 168 7787 224 7789
rect 421 7841 477 7843
rect 421 7789 423 7841
rect 423 7789 475 7841
rect 475 7789 477 7841
rect 421 7787 477 7789
rect 789 7841 845 7843
rect 789 7789 791 7841
rect 791 7789 843 7841
rect 843 7789 845 7841
rect 789 7787 845 7789
rect 1157 7841 1213 7843
rect 1157 7789 1159 7841
rect 1159 7789 1211 7841
rect 1211 7789 1213 7841
rect 1157 7787 1213 7789
rect 1525 7841 1581 7843
rect 1525 7789 1527 7841
rect 1527 7789 1579 7841
rect 1579 7789 1581 7841
rect 1525 7787 1581 7789
rect 628 7096 684 7098
rect 628 7044 630 7096
rect 630 7044 682 7096
rect 682 7044 684 7096
rect 628 7042 684 7044
rect 1364 7096 1420 7098
rect 1364 7044 1366 7096
rect 1366 7044 1418 7096
rect 1418 7044 1420 7096
rect 1364 7042 1420 7044
rect 168 6351 224 6353
rect 168 6299 170 6351
rect 170 6299 222 6351
rect 222 6299 224 6351
rect 168 6297 224 6299
rect 421 6351 477 6353
rect 421 6299 423 6351
rect 423 6299 475 6351
rect 475 6299 477 6351
rect 421 6297 477 6299
rect 789 6351 845 6353
rect 789 6299 791 6351
rect 791 6299 843 6351
rect 843 6299 845 6351
rect 789 6297 845 6299
rect 1157 6351 1213 6353
rect 1157 6299 1159 6351
rect 1159 6299 1211 6351
rect 1211 6299 1213 6351
rect 1157 6297 1213 6299
rect 1525 6351 1581 6353
rect 1525 6299 1527 6351
rect 1527 6299 1579 6351
rect 1579 6299 1581 6351
rect 1525 6297 1581 6299
rect 628 5682 684 5684
rect 628 5630 630 5682
rect 630 5630 682 5682
rect 682 5630 684 5682
rect 628 5628 684 5630
rect 1364 5682 1420 5684
rect 1364 5630 1366 5682
rect 1366 5630 1418 5682
rect 1418 5630 1420 5682
rect 1364 5628 1420 5630
rect 168 5013 224 5015
rect 168 4961 170 5013
rect 170 4961 222 5013
rect 222 4961 224 5013
rect 168 4959 224 4961
rect 421 5013 477 5015
rect 421 4961 423 5013
rect 423 4961 475 5013
rect 475 4961 477 5013
rect 421 4959 477 4961
rect 789 5013 845 5015
rect 789 4961 791 5013
rect 791 4961 843 5013
rect 843 4961 845 5013
rect 789 4959 845 4961
rect 1157 5013 1213 5015
rect 1157 4961 1159 5013
rect 1159 4961 1211 5013
rect 1211 4961 1213 5013
rect 1157 4959 1213 4961
rect 1525 5013 1581 5015
rect 1525 4961 1527 5013
rect 1527 4961 1579 5013
rect 1579 4961 1581 5013
rect 1525 4959 1581 4961
rect 628 4268 684 4270
rect 628 4216 630 4268
rect 630 4216 682 4268
rect 682 4216 684 4268
rect 628 4214 684 4216
rect 1364 4268 1420 4270
rect 1364 4216 1366 4268
rect 1366 4216 1418 4268
rect 1418 4216 1420 4268
rect 1364 4214 1420 4216
rect 168 3523 224 3525
rect 168 3471 170 3523
rect 170 3471 222 3523
rect 222 3471 224 3523
rect 168 3469 224 3471
rect 421 3523 477 3525
rect 421 3471 423 3523
rect 423 3471 475 3523
rect 475 3471 477 3523
rect 421 3469 477 3471
rect 789 3523 845 3525
rect 789 3471 791 3523
rect 791 3471 843 3523
rect 843 3471 845 3523
rect 789 3469 845 3471
rect 1157 3523 1213 3525
rect 1157 3471 1159 3523
rect 1159 3471 1211 3523
rect 1211 3471 1213 3523
rect 1157 3469 1213 3471
rect 1525 3523 1581 3525
rect 1525 3471 1527 3523
rect 1527 3471 1579 3523
rect 1579 3471 1581 3523
rect 1525 3469 1581 3471
rect 628 2854 684 2856
rect 628 2802 630 2854
rect 630 2802 682 2854
rect 682 2802 684 2854
rect 628 2800 684 2802
rect 1364 2854 1420 2856
rect 1364 2802 1366 2854
rect 1366 2802 1418 2854
rect 1418 2802 1420 2854
rect 1364 2800 1420 2802
rect 168 2185 224 2187
rect 168 2133 170 2185
rect 170 2133 222 2185
rect 222 2133 224 2185
rect 168 2131 224 2133
rect 421 2185 477 2187
rect 421 2133 423 2185
rect 423 2133 475 2185
rect 475 2133 477 2185
rect 421 2131 477 2133
rect 789 2185 845 2187
rect 789 2133 791 2185
rect 791 2133 843 2185
rect 843 2133 845 2185
rect 789 2131 845 2133
rect 1157 2185 1213 2187
rect 1157 2133 1159 2185
rect 1159 2133 1211 2185
rect 1211 2133 1213 2185
rect 1157 2131 1213 2133
rect 1525 2185 1581 2187
rect 1525 2133 1527 2185
rect 1527 2133 1579 2185
rect 1579 2133 1581 2185
rect 1525 2131 1581 2133
rect 628 1440 684 1442
rect 628 1388 630 1440
rect 630 1388 682 1440
rect 682 1388 684 1440
rect 628 1386 684 1388
rect 1364 1440 1420 1442
rect 1364 1388 1366 1440
rect 1366 1388 1418 1440
rect 1418 1388 1420 1440
rect 1364 1386 1420 1388
rect 168 695 224 697
rect 168 643 170 695
rect 170 643 222 695
rect 222 643 224 695
rect 168 641 224 643
rect 421 695 477 697
rect 421 643 423 695
rect 423 643 475 695
rect 475 643 477 695
rect 421 641 477 643
rect 789 695 845 697
rect 789 643 791 695
rect 791 643 843 695
rect 843 643 845 695
rect 789 641 845 643
rect 1157 695 1213 697
rect 1157 643 1159 695
rect 1159 643 1211 695
rect 1211 643 1213 695
rect 1157 641 1213 643
rect 1525 695 1581 697
rect 1525 643 1527 695
rect 1527 643 1579 695
rect 1579 643 1581 695
rect 1525 641 1581 643
rect 628 26 684 28
rect 628 -26 630 26
rect 630 -26 682 26
rect 682 -26 684 26
rect 628 -28 684 -26
rect 1364 26 1420 28
rect 1364 -26 1366 26
rect 1366 -26 1418 26
rect 1418 -26 1420 26
rect 1364 -28 1420 -26
<< metal3 >>
rect 607 12754 705 12775
rect 607 12698 628 12754
rect 684 12698 705 12754
rect 607 12677 705 12698
rect 1343 12754 1441 12775
rect 1343 12698 1364 12754
rect 1420 12698 1441 12754
rect 1343 12677 1441 12698
rect 163 12011 229 12014
rect 416 12011 482 12014
rect 784 12011 850 12014
rect 1152 12011 1218 12014
rect 1520 12011 1586 12014
rect 163 12009 1586 12011
rect 163 11953 168 12009
rect 224 11953 421 12009
rect 477 11953 789 12009
rect 845 11953 1157 12009
rect 1213 11953 1525 12009
rect 1581 11953 1586 12009
rect 163 11951 1586 11953
rect 163 11948 229 11951
rect 416 11948 482 11951
rect 784 11948 850 11951
rect 1152 11948 1218 11951
rect 1520 11948 1586 11951
rect 607 11340 705 11361
rect 607 11284 628 11340
rect 684 11284 705 11340
rect 607 11263 705 11284
rect 1343 11340 1441 11361
rect 1343 11284 1364 11340
rect 1420 11284 1441 11340
rect 1343 11263 1441 11284
rect 163 10673 229 10676
rect 416 10673 482 10676
rect 784 10673 850 10676
rect 1152 10673 1218 10676
rect 1520 10673 1586 10676
rect 163 10671 1586 10673
rect 163 10615 168 10671
rect 224 10615 421 10671
rect 477 10615 789 10671
rect 845 10615 1157 10671
rect 1213 10615 1525 10671
rect 1581 10615 1586 10671
rect 163 10613 1586 10615
rect 163 10610 229 10613
rect 416 10610 482 10613
rect 784 10610 850 10613
rect 1152 10610 1218 10613
rect 1520 10610 1586 10613
rect 607 9926 705 9947
rect 607 9870 628 9926
rect 684 9870 705 9926
rect 607 9849 705 9870
rect 1343 9926 1441 9947
rect 1343 9870 1364 9926
rect 1420 9870 1441 9926
rect 1343 9849 1441 9870
rect 163 9183 229 9186
rect 416 9183 482 9186
rect 784 9183 850 9186
rect 1152 9183 1218 9186
rect 1520 9183 1586 9186
rect 163 9181 1586 9183
rect 163 9125 168 9181
rect 224 9125 421 9181
rect 477 9125 789 9181
rect 845 9125 1157 9181
rect 1213 9125 1525 9181
rect 1581 9125 1586 9181
rect 163 9123 1586 9125
rect 163 9120 229 9123
rect 416 9120 482 9123
rect 784 9120 850 9123
rect 1152 9120 1218 9123
rect 1520 9120 1586 9123
rect 607 8512 705 8533
rect 607 8456 628 8512
rect 684 8456 705 8512
rect 607 8435 705 8456
rect 1343 8512 1441 8533
rect 1343 8456 1364 8512
rect 1420 8456 1441 8512
rect 1343 8435 1441 8456
rect 163 7845 229 7848
rect 416 7845 482 7848
rect 784 7845 850 7848
rect 1152 7845 1218 7848
rect 1520 7845 1586 7848
rect 163 7843 1586 7845
rect 163 7787 168 7843
rect 224 7787 421 7843
rect 477 7787 789 7843
rect 845 7787 1157 7843
rect 1213 7787 1525 7843
rect 1581 7787 1586 7843
rect 163 7785 1586 7787
rect 163 7782 229 7785
rect 416 7782 482 7785
rect 784 7782 850 7785
rect 1152 7782 1218 7785
rect 1520 7782 1586 7785
rect 607 7098 705 7119
rect 607 7042 628 7098
rect 684 7042 705 7098
rect 607 7021 705 7042
rect 1343 7098 1441 7119
rect 1343 7042 1364 7098
rect 1420 7042 1441 7098
rect 1343 7021 1441 7042
rect 163 6355 229 6358
rect 416 6355 482 6358
rect 784 6355 850 6358
rect 1152 6355 1218 6358
rect 1520 6355 1586 6358
rect 163 6353 1586 6355
rect 163 6297 168 6353
rect 224 6297 421 6353
rect 477 6297 789 6353
rect 845 6297 1157 6353
rect 1213 6297 1525 6353
rect 1581 6297 1586 6353
rect 163 6295 1586 6297
rect 163 6292 229 6295
rect 416 6292 482 6295
rect 784 6292 850 6295
rect 1152 6292 1218 6295
rect 1520 6292 1586 6295
rect 607 5684 705 5705
rect 607 5628 628 5684
rect 684 5628 705 5684
rect 607 5607 705 5628
rect 1343 5684 1441 5705
rect 1343 5628 1364 5684
rect 1420 5628 1441 5684
rect 1343 5607 1441 5628
rect 163 5017 229 5020
rect 416 5017 482 5020
rect 784 5017 850 5020
rect 1152 5017 1218 5020
rect 1520 5017 1586 5020
rect 163 5015 1586 5017
rect 163 4959 168 5015
rect 224 4959 421 5015
rect 477 4959 789 5015
rect 845 4959 1157 5015
rect 1213 4959 1525 5015
rect 1581 4959 1586 5015
rect 163 4957 1586 4959
rect 163 4954 229 4957
rect 416 4954 482 4957
rect 784 4954 850 4957
rect 1152 4954 1218 4957
rect 1520 4954 1586 4957
rect 607 4270 705 4291
rect 607 4214 628 4270
rect 684 4214 705 4270
rect 607 4193 705 4214
rect 1343 4270 1441 4291
rect 1343 4214 1364 4270
rect 1420 4214 1441 4270
rect 1343 4193 1441 4214
rect 163 3527 229 3530
rect 416 3527 482 3530
rect 784 3527 850 3530
rect 1152 3527 1218 3530
rect 1520 3527 1586 3530
rect 163 3525 1586 3527
rect 163 3469 168 3525
rect 224 3469 421 3525
rect 477 3469 789 3525
rect 845 3469 1157 3525
rect 1213 3469 1525 3525
rect 1581 3469 1586 3525
rect 163 3467 1586 3469
rect 163 3464 229 3467
rect 416 3464 482 3467
rect 784 3464 850 3467
rect 1152 3464 1218 3467
rect 1520 3464 1586 3467
rect 607 2856 705 2877
rect 607 2800 628 2856
rect 684 2800 705 2856
rect 607 2779 705 2800
rect 1343 2856 1441 2877
rect 1343 2800 1364 2856
rect 1420 2800 1441 2856
rect 1343 2779 1441 2800
rect 163 2189 229 2192
rect 416 2189 482 2192
rect 784 2189 850 2192
rect 1152 2189 1218 2192
rect 1520 2189 1586 2192
rect 163 2187 1586 2189
rect 163 2131 168 2187
rect 224 2131 421 2187
rect 477 2131 789 2187
rect 845 2131 1157 2187
rect 1213 2131 1525 2187
rect 1581 2131 1586 2187
rect 163 2129 1586 2131
rect 163 2126 229 2129
rect 416 2126 482 2129
rect 784 2126 850 2129
rect 1152 2126 1218 2129
rect 1520 2126 1586 2129
rect 607 1442 705 1463
rect 607 1386 628 1442
rect 684 1386 705 1442
rect 607 1365 705 1386
rect 1343 1442 1441 1463
rect 1343 1386 1364 1442
rect 1420 1386 1441 1442
rect 1343 1365 1441 1386
rect 163 699 229 702
rect 416 699 482 702
rect 784 699 850 702
rect 1152 699 1218 702
rect 1520 699 1586 702
rect 163 697 1586 699
rect 163 641 168 697
rect 224 641 421 697
rect 477 641 789 697
rect 845 641 1157 697
rect 1213 641 1525 697
rect 1581 641 1586 697
rect 163 639 1586 641
rect 163 636 229 639
rect 416 636 482 639
rect 784 636 850 639
rect 1152 636 1218 639
rect 1520 636 1586 639
rect 607 28 705 49
rect 607 -28 628 28
rect 684 -28 705 28
rect 607 -49 705 -28
rect 1343 28 1441 49
rect 1343 -28 1364 28
rect 1420 -28 1441 28
rect 1343 -49 1441 -28
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 1524 0 1 11948
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 -75 0 1 637
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 -72 0 1 636
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 1359 0 1 11275
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 1360 0 1 11280
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 1363 0 1 11279
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 623 0 1 11275
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 624 0 1 11280
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 627 0 1 11279
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 1359 0 1 12689
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 1360 0 1 12694
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 1363 0 1 12693
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 623 0 1 12689
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 624 0 1 12694
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 627 0 1 12693
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 1359 0 1 11275
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 1360 0 1 11280
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 1363 0 1 11279
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 623 0 1 11275
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 624 0 1 11280
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 627 0 1 11279
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 1359 0 1 9861
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 1360 0 1 9866
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 1363 0 1 9865
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 623 0 1 9861
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 624 0 1 9866
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 627 0 1 9865
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 1359 0 1 8447
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 1360 0 1 8452
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 1363 0 1 8451
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 623 0 1 8447
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 624 0 1 8452
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 627 0 1 8451
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 1359 0 1 9861
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 1360 0 1 9866
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1634918361
transform 1 0 1363 0 1 9865
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 623 0 1 9861
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 624 0 1 9866
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1634918361
transform 1 0 627 0 1 9865
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 1359 0 1 8447
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 1360 0 1 8452
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1634918361
transform 1 0 1363 0 1 8451
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 623 0 1 8447
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 624 0 1 8452
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1634918361
transform 1 0 627 0 1 8451
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 1359 0 1 7033
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 1360 0 1 7038
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1634918361
transform 1 0 1363 0 1 7037
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 623 0 1 7033
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1634918361
transform 1 0 624 0 1 7038
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1634918361
transform 1 0 627 0 1 7037
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 1359 0 1 5619
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1634918361
transform 1 0 1360 0 1 5624
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1634918361
transform 1 0 1363 0 1 5623
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1634918361
transform 1 0 623 0 1 5619
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1634918361
transform 1 0 624 0 1 5624
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1634918361
transform 1 0 627 0 1 5623
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1634918361
transform 1 0 1359 0 1 7033
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1634918361
transform 1 0 1360 0 1 7038
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1634918361
transform 1 0 1363 0 1 7037
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1634918361
transform 1 0 623 0 1 7033
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1634918361
transform 1 0 624 0 1 7038
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1634918361
transform 1 0 627 0 1 7037
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1634918361
transform 1 0 1359 0 1 5619
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1634918361
transform 1 0 1360 0 1 5624
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1634918361
transform 1 0 1363 0 1 5623
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1634918361
transform 1 0 623 0 1 5619
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1634918361
transform 1 0 624 0 1 5624
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1634918361
transform 1 0 627 0 1 5623
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1634918361
transform 1 0 1359 0 1 4205
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1634918361
transform 1 0 1360 0 1 4210
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1634918361
transform 1 0 1363 0 1 4209
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1634918361
transform 1 0 623 0 1 4205
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1634918361
transform 1 0 624 0 1 4210
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1634918361
transform 1 0 627 0 1 4209
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1634918361
transform 1 0 1359 0 1 2791
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1634918361
transform 1 0 1360 0 1 2796
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1634918361
transform 1 0 1363 0 1 2795
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1634918361
transform 1 0 623 0 1 2791
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1634918361
transform 1 0 624 0 1 2796
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1634918361
transform 1 0 627 0 1 2795
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1634918361
transform 1 0 1359 0 1 4205
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1634918361
transform 1 0 1360 0 1 4210
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1634918361
transform 1 0 1363 0 1 4209
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1634918361
transform 1 0 623 0 1 4205
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1634918361
transform 1 0 624 0 1 4210
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1634918361
transform 1 0 627 0 1 4209
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1634918361
transform 1 0 1359 0 1 2791
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1634918361
transform 1 0 1360 0 1 2796
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1634918361
transform 1 0 1363 0 1 2795
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1634918361
transform 1 0 623 0 1 2791
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1634918361
transform 1 0 624 0 1 2796
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1634918361
transform 1 0 627 0 1 2795
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1634918361
transform 1 0 1359 0 1 1377
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1634918361
transform 1 0 1360 0 1 1382
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1634918361
transform 1 0 1363 0 1 1381
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1634918361
transform 1 0 623 0 1 1377
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1634918361
transform 1 0 624 0 1 1382
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1634918361
transform 1 0 627 0 1 1381
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1634918361
transform 1 0 1359 0 1 -37
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1634918361
transform 1 0 1360 0 1 -32
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1634918361
transform 1 0 1363 0 1 -33
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1634918361
transform 1 0 623 0 1 -37
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1634918361
transform 1 0 624 0 1 -32
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1634918361
transform 1 0 627 0 1 -33
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1634918361
transform 1 0 1359 0 1 1377
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1634918361
transform 1 0 1360 0 1 1382
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1634918361
transform 1 0 1363 0 1 1381
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1634918361
transform 1 0 623 0 1 1377
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1634918361
transform 1 0 624 0 1 1382
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1634918361
transform 1 0 627 0 1 1381
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1634918361
transform 1 0 163 0 1 11944
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1634918361
transform 1 0 164 0 1 11949
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1634918361
transform 1 0 167 0 1 11948
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1634918361
transform 1 0 49 0 1 11949
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1634918361
transform 1 0 52 0 1 11948
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1634918361
transform 1 0 1520 0 1 11944
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1634918361
transform 1 0 1521 0 1 11949
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1634918361
transform 1 0 1524 0 1 11948
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1634918361
transform 1 0 1152 0 1 11944
box 0 0 1 1
use contact_19  contact_19_40
timestamp 1634918361
transform 1 0 1153 0 1 11949
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1634918361
transform 1 0 1156 0 1 11948
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1634918361
transform 1 0 784 0 1 11944
box 0 0 1 1
use contact_19  contact_19_41
timestamp 1634918361
transform 1 0 785 0 1 11949
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1634918361
transform 1 0 788 0 1 11948
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1634918361
transform 1 0 416 0 1 11944
box 0 0 1 1
use contact_19  contact_19_42
timestamp 1634918361
transform 1 0 417 0 1 11949
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1634918361
transform 1 0 420 0 1 11948
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1634918361
transform 1 0 163 0 1 10606
box 0 0 1 1
use contact_19  contact_19_43
timestamp 1634918361
transform 1 0 164 0 1 10611
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1634918361
transform 1 0 167 0 1 10610
box 0 0 1 1
use contact_19  contact_19_44
timestamp 1634918361
transform 1 0 49 0 1 10611
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1634918361
transform 1 0 52 0 1 10610
box 0 0 1 1
use contact_7  contact_7_42
timestamp 1634918361
transform 1 0 1520 0 1 10606
box 0 0 1 1
use contact_19  contact_19_45
timestamp 1634918361
transform 1 0 1521 0 1 10611
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1634918361
transform 1 0 1524 0 1 10610
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1634918361
transform 1 0 1152 0 1 10606
box 0 0 1 1
use contact_19  contact_19_46
timestamp 1634918361
transform 1 0 1153 0 1 10611
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1634918361
transform 1 0 1156 0 1 10610
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1634918361
transform 1 0 784 0 1 10606
box 0 0 1 1
use contact_19  contact_19_47
timestamp 1634918361
transform 1 0 785 0 1 10611
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1634918361
transform 1 0 788 0 1 10610
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1634918361
transform 1 0 416 0 1 10606
box 0 0 1 1
use contact_19  contact_19_48
timestamp 1634918361
transform 1 0 417 0 1 10611
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1634918361
transform 1 0 420 0 1 10610
box 0 0 1 1
use contact_7  contact_7_46
timestamp 1634918361
transform 1 0 163 0 1 9116
box 0 0 1 1
use contact_19  contact_19_49
timestamp 1634918361
transform 1 0 164 0 1 9121
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1634918361
transform 1 0 167 0 1 9120
box 0 0 1 1
use contact_19  contact_19_50
timestamp 1634918361
transform 1 0 49 0 1 9121
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1634918361
transform 1 0 52 0 1 9120
box 0 0 1 1
use contact_7  contact_7_47
timestamp 1634918361
transform 1 0 1520 0 1 9116
box 0 0 1 1
use contact_19  contact_19_51
timestamp 1634918361
transform 1 0 1521 0 1 9121
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1634918361
transform 1 0 1524 0 1 9120
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1634918361
transform 1 0 1152 0 1 9116
box 0 0 1 1
use contact_19  contact_19_52
timestamp 1634918361
transform 1 0 1153 0 1 9121
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1634918361
transform 1 0 1156 0 1 9120
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1634918361
transform 1 0 784 0 1 9116
box 0 0 1 1
use contact_19  contact_19_53
timestamp 1634918361
transform 1 0 785 0 1 9121
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1634918361
transform 1 0 788 0 1 9120
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1634918361
transform 1 0 416 0 1 9116
box 0 0 1 1
use contact_19  contact_19_54
timestamp 1634918361
transform 1 0 417 0 1 9121
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1634918361
transform 1 0 420 0 1 9120
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1634918361
transform 1 0 163 0 1 7778
box 0 0 1 1
use contact_19  contact_19_55
timestamp 1634918361
transform 1 0 164 0 1 7783
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1634918361
transform 1 0 167 0 1 7782
box 0 0 1 1
use contact_19  contact_19_56
timestamp 1634918361
transform 1 0 49 0 1 7783
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1634918361
transform 1 0 52 0 1 7782
box 0 0 1 1
use contact_7  contact_7_52
timestamp 1634918361
transform 1 0 1520 0 1 7778
box 0 0 1 1
use contact_19  contact_19_57
timestamp 1634918361
transform 1 0 1521 0 1 7783
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1634918361
transform 1 0 1524 0 1 7782
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1634918361
transform 1 0 1152 0 1 7778
box 0 0 1 1
use contact_19  contact_19_58
timestamp 1634918361
transform 1 0 1153 0 1 7783
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1634918361
transform 1 0 1156 0 1 7782
box 0 0 1 1
use contact_7  contact_7_54
timestamp 1634918361
transform 1 0 784 0 1 7778
box 0 0 1 1
use contact_19  contact_19_59
timestamp 1634918361
transform 1 0 785 0 1 7783
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1634918361
transform 1 0 788 0 1 7782
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1634918361
transform 1 0 416 0 1 7778
box 0 0 1 1
use contact_19  contact_19_60
timestamp 1634918361
transform 1 0 417 0 1 7783
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1634918361
transform 1 0 420 0 1 7782
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1634918361
transform 1 0 163 0 1 6288
box 0 0 1 1
use contact_19  contact_19_61
timestamp 1634918361
transform 1 0 164 0 1 6293
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1634918361
transform 1 0 167 0 1 6292
box 0 0 1 1
use contact_19  contact_19_62
timestamp 1634918361
transform 1 0 49 0 1 6293
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1634918361
transform 1 0 52 0 1 6292
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1634918361
transform 1 0 1520 0 1 6288
box 0 0 1 1
use contact_19  contact_19_63
timestamp 1634918361
transform 1 0 1521 0 1 6293
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1634918361
transform 1 0 1524 0 1 6292
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1634918361
transform 1 0 1152 0 1 6288
box 0 0 1 1
use contact_19  contact_19_64
timestamp 1634918361
transform 1 0 1153 0 1 6293
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1634918361
transform 1 0 1156 0 1 6292
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1634918361
transform 1 0 784 0 1 6288
box 0 0 1 1
use contact_19  contact_19_65
timestamp 1634918361
transform 1 0 785 0 1 6293
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1634918361
transform 1 0 788 0 1 6292
box 0 0 1 1
use contact_7  contact_7_60
timestamp 1634918361
transform 1 0 416 0 1 6288
box 0 0 1 1
use contact_19  contact_19_66
timestamp 1634918361
transform 1 0 417 0 1 6293
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1634918361
transform 1 0 420 0 1 6292
box 0 0 1 1
use contact_7  contact_7_61
timestamp 1634918361
transform 1 0 163 0 1 4950
box 0 0 1 1
use contact_19  contact_19_67
timestamp 1634918361
transform 1 0 164 0 1 4955
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1634918361
transform 1 0 167 0 1 4954
box 0 0 1 1
use contact_19  contact_19_68
timestamp 1634918361
transform 1 0 49 0 1 4955
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1634918361
transform 1 0 52 0 1 4954
box 0 0 1 1
use contact_7  contact_7_62
timestamp 1634918361
transform 1 0 1520 0 1 4950
box 0 0 1 1
use contact_19  contact_19_69
timestamp 1634918361
transform 1 0 1521 0 1 4955
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1634918361
transform 1 0 1524 0 1 4954
box 0 0 1 1
use contact_7  contact_7_63
timestamp 1634918361
transform 1 0 1152 0 1 4950
box 0 0 1 1
use contact_19  contact_19_70
timestamp 1634918361
transform 1 0 1153 0 1 4955
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1634918361
transform 1 0 1156 0 1 4954
box 0 0 1 1
use contact_7  contact_7_64
timestamp 1634918361
transform 1 0 784 0 1 4950
box 0 0 1 1
use contact_19  contact_19_71
timestamp 1634918361
transform 1 0 785 0 1 4955
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1634918361
transform 1 0 788 0 1 4954
box 0 0 1 1
use contact_7  contact_7_65
timestamp 1634918361
transform 1 0 416 0 1 4950
box 0 0 1 1
use contact_19  contact_19_72
timestamp 1634918361
transform 1 0 417 0 1 4955
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1634918361
transform 1 0 420 0 1 4954
box 0 0 1 1
use contact_7  contact_7_66
timestamp 1634918361
transform 1 0 163 0 1 3460
box 0 0 1 1
use contact_19  contact_19_73
timestamp 1634918361
transform 1 0 164 0 1 3465
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1634918361
transform 1 0 167 0 1 3464
box 0 0 1 1
use contact_19  contact_19_74
timestamp 1634918361
transform 1 0 49 0 1 3465
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1634918361
transform 1 0 52 0 1 3464
box 0 0 1 1
use contact_7  contact_7_67
timestamp 1634918361
transform 1 0 1520 0 1 3460
box 0 0 1 1
use contact_19  contact_19_75
timestamp 1634918361
transform 1 0 1521 0 1 3465
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1634918361
transform 1 0 1524 0 1 3464
box 0 0 1 1
use contact_7  contact_7_68
timestamp 1634918361
transform 1 0 1152 0 1 3460
box 0 0 1 1
use contact_19  contact_19_76
timestamp 1634918361
transform 1 0 1153 0 1 3465
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1634918361
transform 1 0 1156 0 1 3464
box 0 0 1 1
use contact_7  contact_7_69
timestamp 1634918361
transform 1 0 784 0 1 3460
box 0 0 1 1
use contact_19  contact_19_77
timestamp 1634918361
transform 1 0 785 0 1 3465
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1634918361
transform 1 0 788 0 1 3464
box 0 0 1 1
use contact_7  contact_7_70
timestamp 1634918361
transform 1 0 416 0 1 3460
box 0 0 1 1
use contact_19  contact_19_78
timestamp 1634918361
transform 1 0 417 0 1 3465
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1634918361
transform 1 0 420 0 1 3464
box 0 0 1 1
use contact_7  contact_7_71
timestamp 1634918361
transform 1 0 163 0 1 2122
box 0 0 1 1
use contact_19  contact_19_79
timestamp 1634918361
transform 1 0 164 0 1 2127
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1634918361
transform 1 0 167 0 1 2126
box 0 0 1 1
use contact_19  contact_19_80
timestamp 1634918361
transform 1 0 49 0 1 2127
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1634918361
transform 1 0 52 0 1 2126
box 0 0 1 1
use contact_7  contact_7_72
timestamp 1634918361
transform 1 0 1520 0 1 2122
box 0 0 1 1
use contact_19  contact_19_81
timestamp 1634918361
transform 1 0 1521 0 1 2127
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1634918361
transform 1 0 1524 0 1 2126
box 0 0 1 1
use contact_7  contact_7_73
timestamp 1634918361
transform 1 0 1152 0 1 2122
box 0 0 1 1
use contact_19  contact_19_82
timestamp 1634918361
transform 1 0 1153 0 1 2127
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1634918361
transform 1 0 1156 0 1 2126
box 0 0 1 1
use contact_7  contact_7_74
timestamp 1634918361
transform 1 0 784 0 1 2122
box 0 0 1 1
use contact_19  contact_19_83
timestamp 1634918361
transform 1 0 785 0 1 2127
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1634918361
transform 1 0 788 0 1 2126
box 0 0 1 1
use contact_7  contact_7_75
timestamp 1634918361
transform 1 0 416 0 1 2122
box 0 0 1 1
use contact_19  contact_19_84
timestamp 1634918361
transform 1 0 417 0 1 2127
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1634918361
transform 1 0 420 0 1 2126
box 0 0 1 1
use contact_7  contact_7_76
timestamp 1634918361
transform 1 0 163 0 1 632
box 0 0 1 1
use contact_19  contact_19_85
timestamp 1634918361
transform 1 0 164 0 1 637
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1634918361
transform 1 0 167 0 1 636
box 0 0 1 1
use contact_19  contact_19_86
timestamp 1634918361
transform 1 0 49 0 1 637
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1634918361
transform 1 0 52 0 1 636
box 0 0 1 1
use contact_7  contact_7_77
timestamp 1634918361
transform 1 0 1520 0 1 632
box 0 0 1 1
use contact_19  contact_19_87
timestamp 1634918361
transform 1 0 1521 0 1 637
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1634918361
transform 1 0 1524 0 1 636
box 0 0 1 1
use contact_7  contact_7_78
timestamp 1634918361
transform 1 0 1152 0 1 632
box 0 0 1 1
use contact_19  contact_19_88
timestamp 1634918361
transform 1 0 1153 0 1 637
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1634918361
transform 1 0 1156 0 1 636
box 0 0 1 1
use contact_7  contact_7_79
timestamp 1634918361
transform 1 0 784 0 1 632
box 0 0 1 1
use contact_19  contact_19_89
timestamp 1634918361
transform 1 0 785 0 1 637
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1634918361
transform 1 0 788 0 1 636
box 0 0 1 1
use contact_7  contact_7_80
timestamp 1634918361
transform 1 0 416 0 1 632
box 0 0 1 1
use contact_19  contact_19_90
timestamp 1634918361
transform 1 0 417 0 1 637
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1634918361
transform 1 0 420 0 1 636
box 0 0 1 1
use pinv_11  pinv_11_0
timestamp 1634918361
transform 1 0 1472 0 1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_1
timestamp 1634918361
transform 1 0 1104 0 1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_2
timestamp 1634918361
transform 1 0 736 0 1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_3
timestamp 1634918361
transform 1 0 368 0 1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_4
timestamp 1634918361
transform 1 0 0 0 1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_5
timestamp 1634918361
transform 1 0 1472 0 -1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_6
timestamp 1634918361
transform 1 0 1104 0 -1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_7
timestamp 1634918361
transform 1 0 736 0 -1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_8
timestamp 1634918361
transform 1 0 368 0 -1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_9
timestamp 1634918361
transform 1 0 0 0 -1 11312
box -36 -17 404 1471
use pinv_11  pinv_11_10
timestamp 1634918361
transform 1 0 1472 0 1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_11
timestamp 1634918361
transform 1 0 1104 0 1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_12
timestamp 1634918361
transform 1 0 736 0 1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_13
timestamp 1634918361
transform 1 0 368 0 1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_14
timestamp 1634918361
transform 1 0 0 0 1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_15
timestamp 1634918361
transform 1 0 1472 0 -1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_16
timestamp 1634918361
transform 1 0 1104 0 -1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_17
timestamp 1634918361
transform 1 0 736 0 -1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_18
timestamp 1634918361
transform 1 0 368 0 -1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_19
timestamp 1634918361
transform 1 0 0 0 -1 8484
box -36 -17 404 1471
use pinv_11  pinv_11_20
timestamp 1634918361
transform 1 0 1472 0 1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_21
timestamp 1634918361
transform 1 0 1104 0 1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_22
timestamp 1634918361
transform 1 0 736 0 1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_23
timestamp 1634918361
transform 1 0 368 0 1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_24
timestamp 1634918361
transform 1 0 0 0 1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_25
timestamp 1634918361
transform 1 0 1472 0 -1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_26
timestamp 1634918361
transform 1 0 1104 0 -1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_27
timestamp 1634918361
transform 1 0 736 0 -1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_28
timestamp 1634918361
transform 1 0 368 0 -1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_29
timestamp 1634918361
transform 1 0 0 0 -1 5656
box -36 -17 404 1471
use pinv_11  pinv_11_30
timestamp 1634918361
transform 1 0 1472 0 1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_31
timestamp 1634918361
transform 1 0 1104 0 1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_32
timestamp 1634918361
transform 1 0 736 0 1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_33
timestamp 1634918361
transform 1 0 368 0 1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_34
timestamp 1634918361
transform 1 0 0 0 1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_35
timestamp 1634918361
transform 1 0 1472 0 -1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_36
timestamp 1634918361
transform 1 0 1104 0 -1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_37
timestamp 1634918361
transform 1 0 736 0 -1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_38
timestamp 1634918361
transform 1 0 368 0 -1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_39
timestamp 1634918361
transform 1 0 0 0 -1 2828
box -36 -17 404 1471
use pinv_11  pinv_11_40
timestamp 1634918361
transform 1 0 1472 0 1 0
box -36 -17 404 1471
use pinv_11  pinv_11_41
timestamp 1634918361
transform 1 0 1104 0 1 0
box -36 -17 404 1471
use pinv_11  pinv_11_42
timestamp 1634918361
transform 1 0 736 0 1 0
box -36 -17 404 1471
use pinv_11  pinv_11_43
timestamp 1634918361
transform 1 0 368 0 1 0
box -36 -17 404 1471
use pinv_11  pinv_11_44
timestamp 1634918361
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel metal3 s 1343 9849 1441 9947 4 vdd
port 1 nsew
rlabel metal3 s 607 7021 705 7119 4 vdd
port 1 nsew
rlabel metal3 s 1343 1365 1441 1463 4 vdd
port 1 nsew
rlabel metal3 s 607 9849 705 9947 4 vdd
port 1 nsew
rlabel metal3 s 1343 4193 1441 4291 4 vdd
port 1 nsew
rlabel metal3 s 1343 12677 1441 12775 4 vdd
port 1 nsew
rlabel metal3 s 607 1365 705 1463 4 vdd
port 1 nsew
rlabel metal3 s 607 12677 705 12775 4 vdd
port 1 nsew
rlabel metal3 s 1343 7021 1441 7119 4 vdd
port 1 nsew
rlabel metal3 s 607 4193 705 4291 4 vdd
port 1 nsew
rlabel metal3 s 607 2779 705 2877 4 gnd
port 2 nsew
rlabel metal3 s 1343 2779 1441 2877 4 gnd
port 2 nsew
rlabel metal3 s 1343 5607 1441 5705 4 gnd
port 2 nsew
rlabel metal3 s 1343 11263 1441 11361 4 gnd
port 2 nsew
rlabel metal3 s 607 -49 705 49 4 gnd
port 2 nsew
rlabel metal3 s 607 8435 705 8533 4 gnd
port 2 nsew
rlabel metal3 s 607 11263 705 11361 4 gnd
port 2 nsew
rlabel metal3 s 607 5607 705 5705 4 gnd
port 2 nsew
rlabel metal3 s 1343 -49 1441 49 4 gnd
port 2 nsew
rlabel metal3 s 1343 8435 1441 8533 4 gnd
port 2 nsew
rlabel metal2 s -57 655 -29 683 4 in
port 3 nsew
rlabel metal1 s 1539 11967 1567 11995 4 out
port 4 nsew
<< properties >>
string FIXED_BBOX 1359 -37 1425 0
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1172004
string GDS_START 1141568
<< end >>
