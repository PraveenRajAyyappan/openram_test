magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1309 -1309 7675 2437
<< locali >>
rect -17 1137 17 1153
rect -17 1087 17 1103
rect 1730 1137 1764 1153
rect 1730 1087 1764 1103
rect 2978 1137 3012 1153
rect 2978 1087 3012 1103
rect 4226 1137 4260 1153
rect 4226 1087 4260 1103
rect 5474 1137 5508 1153
rect 5474 1087 5508 1103
rect 6349 1137 6383 1153
rect 6349 1087 6383 1103
rect 1586 535 1620 551
rect 1931 505 1965 539
rect 2834 535 2868 551
rect 1586 485 1620 501
rect 3179 505 3213 539
rect 4082 535 4116 551
rect 2834 485 2868 501
rect 4427 505 4461 539
rect 5330 535 5364 551
rect 4082 485 4116 501
rect 5675 505 5709 539
rect 5330 485 5364 501
rect 1357 287 1391 303
rect 2605 287 2639 303
rect 3853 287 3887 303
rect 5101 287 5135 303
rect 1391 253 1503 287
rect 2639 253 2751 287
rect 3887 253 3999 287
rect 5135 253 5247 287
rect 1357 237 1391 253
rect 2605 237 2639 253
rect 3853 237 3887 253
rect 5101 237 5135 253
rect -17 17 17 33
rect -17 -33 17 -17
rect 1730 17 1764 33
rect 1730 -33 1764 -17
rect 2978 17 3012 33
rect 2978 -33 3012 -17
rect 4226 17 4260 33
rect 4226 -33 4260 -17
rect 5474 17 5508 33
rect 5474 -33 5508 -17
rect 6349 17 6383 33
rect 6349 -33 6383 -17
<< viali >>
rect -17 1103 17 1137
rect 1730 1103 1764 1137
rect 2978 1103 3012 1137
rect 4226 1103 4260 1137
rect 5474 1103 5508 1137
rect 6349 1103 6383 1137
rect 1586 501 1620 535
rect 2834 501 2868 535
rect 4082 501 4116 535
rect 5330 501 5364 535
rect 1357 253 1391 287
rect 2605 253 2639 287
rect 3853 253 3887 287
rect 5101 253 5135 287
rect -17 -17 17 17
rect 1730 -17 1764 17
rect 2978 -17 3012 17
rect 4226 -17 4260 17
rect 5474 -17 5508 17
rect 6349 -17 6383 17
<< metal1 >>
rect -32 1094 -26 1146
rect 26 1134 32 1146
rect 1718 1137 1776 1143
rect 1718 1134 1730 1137
rect 26 1106 1730 1134
rect 26 1094 32 1106
rect 1718 1103 1730 1106
rect 1764 1134 1776 1137
rect 2966 1137 3024 1143
rect 2966 1134 2978 1137
rect 1764 1106 2978 1134
rect 1764 1103 1776 1106
rect 1718 1097 1776 1103
rect 2966 1103 2978 1106
rect 3012 1134 3024 1137
rect 4214 1137 4272 1143
rect 4214 1134 4226 1137
rect 3012 1106 4226 1134
rect 3012 1103 3024 1106
rect 2966 1097 3024 1103
rect 4214 1103 4226 1106
rect 4260 1134 4272 1137
rect 5462 1137 5520 1143
rect 5462 1134 5474 1137
rect 4260 1106 5474 1134
rect 4260 1103 4272 1106
rect 4214 1097 4272 1103
rect 5462 1103 5474 1106
rect 5508 1134 5520 1137
rect 6334 1134 6340 1146
rect 5508 1106 6340 1134
rect 5508 1103 5520 1106
rect 5462 1097 5520 1103
rect 6334 1094 6340 1106
rect 6392 1094 6398 1146
rect 1571 492 1577 544
rect 1629 492 1635 544
rect 2819 492 2825 544
rect 2877 492 2883 544
rect 4067 492 4073 544
rect 4125 492 4131 544
rect 5315 492 5321 544
rect 5373 492 5379 544
rect 1342 244 1348 296
rect 1400 244 1406 296
rect 2590 244 2596 296
rect 2648 244 2654 296
rect 3838 244 3844 296
rect 3896 244 3902 296
rect 5086 244 5092 296
rect 5144 244 5150 296
rect -32 -26 -26 26
rect 26 14 32 26
rect 1718 17 1776 23
rect 1718 14 1730 17
rect 26 -14 1730 14
rect 26 -26 32 -14
rect 1718 -17 1730 -14
rect 1764 14 1776 17
rect 2966 17 3024 23
rect 2966 14 2978 17
rect 1764 -14 2978 14
rect 1764 -17 1776 -14
rect 1718 -23 1776 -17
rect 2966 -17 2978 -14
rect 3012 14 3024 17
rect 4214 17 4272 23
rect 4214 14 4226 17
rect 3012 -14 4226 14
rect 3012 -17 3024 -14
rect 2966 -23 3024 -17
rect 4214 -17 4226 -14
rect 4260 14 4272 17
rect 5462 17 5520 23
rect 5462 14 5474 17
rect 4260 -14 5474 14
rect 4260 -17 4272 -14
rect 4214 -23 4272 -17
rect 5462 -17 5474 -14
rect 5508 14 5520 17
rect 6334 14 6340 26
rect 5508 -14 6340 14
rect 5508 -17 5520 -14
rect 5462 -23 5520 -17
rect 6334 -26 6340 -14
rect 6392 -26 6398 26
<< via1 >>
rect -26 1137 26 1146
rect -26 1103 -17 1137
rect -17 1103 17 1137
rect 17 1103 26 1137
rect -26 1094 26 1103
rect 6340 1137 6392 1146
rect 6340 1103 6349 1137
rect 6349 1103 6383 1137
rect 6383 1103 6392 1137
rect 6340 1094 6392 1103
rect 1577 535 1629 544
rect 1577 501 1586 535
rect 1586 501 1620 535
rect 1620 501 1629 535
rect 1577 492 1629 501
rect 2825 535 2877 544
rect 2825 501 2834 535
rect 2834 501 2868 535
rect 2868 501 2877 535
rect 2825 492 2877 501
rect 4073 535 4125 544
rect 4073 501 4082 535
rect 4082 501 4116 535
rect 4116 501 4125 535
rect 4073 492 4125 501
rect 5321 535 5373 544
rect 5321 501 5330 535
rect 5330 501 5364 535
rect 5364 501 5373 535
rect 5321 492 5373 501
rect 1348 287 1400 296
rect 1348 253 1357 287
rect 1357 253 1391 287
rect 1391 253 1400 287
rect 1348 244 1400 253
rect 2596 287 2648 296
rect 2596 253 2605 287
rect 2605 253 2639 287
rect 2639 253 2648 287
rect 2596 244 2648 253
rect 3844 287 3896 296
rect 3844 253 3853 287
rect 3853 253 3887 287
rect 3887 253 3896 287
rect 3844 244 3896 253
rect 5092 287 5144 296
rect 5092 253 5101 287
rect 5101 253 5135 287
rect 5135 253 5144 287
rect 5092 244 5144 253
rect -26 17 26 26
rect -26 -17 -17 17
rect -17 -17 17 17
rect 17 -17 26 17
rect -26 -26 26 -17
rect 6340 17 6392 26
rect 6340 -17 6349 17
rect 6349 -17 6383 17
rect 6383 -17 6392 17
rect 6340 -26 6392 -17
<< metal2 >>
rect -28 1148 28 1157
rect -28 1083 28 1092
rect 6338 1148 6394 1157
rect 6338 1083 6394 1092
rect 1575 546 1631 555
rect 1575 481 1631 490
rect 2823 546 2879 555
rect 2823 481 2879 490
rect 4071 546 4127 555
rect 4071 481 4127 490
rect 5319 546 5375 555
rect 5319 481 5375 490
rect 1348 296 1400 302
rect 1348 238 1400 244
rect 2596 296 2648 302
rect 2596 238 2648 244
rect 3844 296 3896 302
rect 3844 238 3896 244
rect 5092 296 5144 302
rect 5092 238 5144 244
rect -28 28 28 37
rect -28 -37 28 -28
rect 6338 28 6394 37
rect 6338 -37 6394 -28
<< via2 >>
rect -28 1146 28 1148
rect -28 1094 -26 1146
rect -26 1094 26 1146
rect 26 1094 28 1146
rect -28 1092 28 1094
rect 6338 1146 6394 1148
rect 6338 1094 6340 1146
rect 6340 1094 6392 1146
rect 6392 1094 6394 1146
rect 6338 1092 6394 1094
rect 1575 544 1631 546
rect 1575 492 1577 544
rect 1577 492 1629 544
rect 1629 492 1631 544
rect 1575 490 1631 492
rect 2823 544 2879 546
rect 2823 492 2825 544
rect 2825 492 2877 544
rect 2877 492 2879 544
rect 2823 490 2879 492
rect 4071 544 4127 546
rect 4071 492 4073 544
rect 4073 492 4125 544
rect 4125 492 4127 544
rect 4071 490 4127 492
rect 5319 544 5375 546
rect 5319 492 5321 544
rect 5321 492 5373 544
rect 5373 492 5375 544
rect 5319 490 5375 492
rect -28 26 28 28
rect -28 -26 -26 26
rect -26 -26 26 26
rect 26 -26 28 26
rect -28 -28 28 -26
rect 6338 26 6394 28
rect 6338 -26 6340 26
rect 6340 -26 6392 26
rect 6392 -26 6394 26
rect 6338 -28 6394 -26
<< metal3 >>
rect -49 1148 49 1169
rect -49 1092 -28 1148
rect 28 1092 49 1148
rect -49 1071 49 1092
rect 6317 1148 6415 1169
rect 6317 1092 6338 1148
rect 6394 1092 6415 1148
rect 6317 1071 6415 1092
rect 1570 548 1636 551
rect 2818 548 2884 551
rect 4066 548 4132 551
rect 5314 548 5380 551
rect 0 546 6366 548
rect 0 490 1575 546
rect 1631 490 2823 546
rect 2879 490 4071 546
rect 4127 490 5319 546
rect 5375 490 6366 546
rect 0 488 6366 490
rect 1570 485 1636 488
rect 2818 485 2884 488
rect 4066 485 4132 488
rect 5314 485 5380 488
rect -49 28 49 49
rect -49 -28 -28 28
rect 28 -28 49 28
rect -49 -49 49 -28
rect 6317 28 6415 49
rect 6317 -28 6338 28
rect 6394 -28 6415 28
rect 6317 -49 6415 -28
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 6333 0 1 1083
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 6334 0 1 1088
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 6337 0 1 1087
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 6337 0 1 1087
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 -33 0 1 1083
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 -32 0 1 1088
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 -29 0 1 1087
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 -29 0 1 1087
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 6333 0 1 -37
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 6334 0 1 -32
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 6337 0 1 -33
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 6337 0 1 -33
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 -33 0 1 -37
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 -32 0 1 -32
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 -29 0 1 -33
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 -29 0 1 -33
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 5462 0 1 1087
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 5462 0 1 -33
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 5314 0 1 481
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 5315 0 1 486
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 5318 0 1 485
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 5086 0 1 238
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 5089 0 1 237
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1634918361
transform 1 0 4214 0 1 1087
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1634918361
transform 1 0 4214 0 1 -33
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 4066 0 1 481
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 4067 0 1 486
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1634918361
transform 1 0 4070 0 1 485
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 3838 0 1 238
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1634918361
transform 1 0 3841 0 1 237
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1634918361
transform 1 0 2966 0 1 1087
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1634918361
transform 1 0 2966 0 1 -33
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 2818 0 1 481
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 2819 0 1 486
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1634918361
transform 1 0 2822 0 1 485
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 2590 0 1 238
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1634918361
transform 1 0 2593 0 1 237
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1634918361
transform 1 0 1718 0 1 1087
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1634918361
transform 1 0 1718 0 1 -33
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 1570 0 1 481
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 1571 0 1 486
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1634918361
transform 1 0 1574 0 1 485
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 1342 0 1 238
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1634918361
transform 1 0 1345 0 1 237
box 0 0 1 1
use pand2  pand2_0
timestamp 1634918361
transform 1 0 5118 0 1 0
box -36 -17 782 1177
use pand2  pand2_1
timestamp 1634918361
transform 1 0 3870 0 1 0
box -36 -17 782 1177
use pand2  pand2_2
timestamp 1634918361
transform 1 0 2622 0 1 0
box -36 -17 782 1177
use pand2  pand2_3
timestamp 1634918361
transform 1 0 1374 0 1 0
box -36 -17 782 1177
<< labels >>
rlabel metal3 s 0 488 6366 548 4 en
port 1 nsew
rlabel metal2 s 1360 256 1388 284 4 wmask_in_0
port 2 nsew
rlabel locali s 1948 522 1948 522 4 wmask_out_0
port 3 nsew
rlabel metal2 s 2608 256 2636 284 4 wmask_in_1
port 4 nsew
rlabel locali s 3196 522 3196 522 4 wmask_out_1
port 5 nsew
rlabel metal2 s 3856 256 3884 284 4 wmask_in_2
port 6 nsew
rlabel locali s 4444 522 4444 522 4 wmask_out_2
port 7 nsew
rlabel metal2 s 5104 256 5132 284 4 wmask_in_3
port 8 nsew
rlabel locali s 5692 522 5692 522 4 wmask_out_3
port 9 nsew
rlabel metal3 s -49 -49 49 49 4 gnd
port 10 nsew
rlabel metal3 s 6317 -49 6415 49 4 gnd
port 10 nsew
rlabel metal3 s 6317 1071 6415 1169 4 vdd
port 11 nsew
rlabel metal3 s -49 1071 49 1169 4 vdd
port 11 nsew
<< properties >>
string FIXED_BBOX 6333 -37 6399 0
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 874242
string GDS_START 868482
<< end >>
