magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1296 -1277 1664 2437
<< nwell >>
rect -36 538 404 1177
<< locali >>
rect 0 1103 368 1137
rect 64 489 98 555
rect 179 505 213 539
rect 0 -17 368 17
use pinv  pinv_0
timestamp 1634918361
transform 1 0 0 0 1 0
box -36 -17 404 1177
<< labels >>
rlabel locali s 196 522 196 522 4 Z
port 1 nsew
rlabel locali s 81 522 81 522 4 A
port 2 nsew
rlabel locali s 184 0 184 0 4 gnd
port 3 nsew
rlabel locali s 184 1120 184 1120 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1120
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 881306
string GDS_START 880512
<< end >>
