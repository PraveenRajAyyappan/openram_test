magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1286 -1286 1868 1652
<< pwell >>
rect -26 -26 608 362
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
rect 384 0 414 336
rect 492 0 522 336
<< ndiff >>
rect 0 185 60 336
rect 0 151 8 185
rect 42 151 60 185
rect 0 0 60 151
rect 90 185 168 336
rect 90 151 112 185
rect 146 151 168 185
rect 90 0 168 151
rect 198 185 276 336
rect 198 151 220 185
rect 254 151 276 185
rect 198 0 276 151
rect 306 185 384 336
rect 306 151 328 185
rect 362 151 384 185
rect 306 0 384 151
rect 414 185 492 336
rect 414 151 436 185
rect 470 151 492 185
rect 414 0 492 151
rect 522 185 582 336
rect 522 151 540 185
rect 574 151 582 185
rect 522 0 582 151
<< ndiffc >>
rect 8 151 42 185
rect 112 151 146 185
rect 220 151 254 185
rect 328 151 362 185
rect 436 151 470 185
rect 540 151 574 185
<< poly >>
rect 60 362 522 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 384 336 414 362
rect 492 336 522 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
<< locali >>
rect 112 235 574 269
rect 8 185 42 201
rect 8 135 42 151
rect 112 185 146 235
rect 112 135 146 151
rect 220 185 254 201
rect 220 135 254 151
rect 328 185 362 235
rect 328 135 362 151
rect 436 185 470 201
rect 436 135 470 151
rect 540 185 574 235
rect 540 135 574 151
use contact_11  contact_11_0
timestamp 1634918361
transform 1 0 532 0 1 135
box 0 0 1 1
use contact_11  contact_11_1
timestamp 1634918361
transform 1 0 428 0 1 135
box 0 0 1 1
use contact_11  contact_11_2
timestamp 1634918361
transform 1 0 320 0 1 135
box 0 0 1 1
use contact_11  contact_11_3
timestamp 1634918361
transform 1 0 212 0 1 135
box 0 0 1 1
use contact_11  contact_11_4
timestamp 1634918361
transform 1 0 104 0 1 135
box 0 0 1 1
use contact_11  contact_11_5
timestamp 1634918361
transform 1 0 0 0 1 135
box 0 0 1 1
<< labels >>
rlabel poly s 291 377 291 377 4 G
port 1 nsew
rlabel locali s 237 168 237 168 4 S
port 2 nsew
rlabel locali s 25 168 25 168 4 S
port 2 nsew
rlabel locali s 453 168 453 168 4 S
port 2 nsew
rlabel locali s 343 252 343 252 4 D
port 3 nsew
<< properties >>
string FIXED_BBOX -25 -26 607 392
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1099836
string GDS_START 1098284
<< end >>
