magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -262 -1256 7878 3271
<< metal1 >>
rect 1500 1959 1530 2011
rect 1702 1959 1732 2011
rect 2140 1959 2170 2011
rect 2342 1959 2372 2011
rect 2748 1959 2778 2011
rect 2950 1959 2980 2011
rect 3388 1959 3418 2011
rect 3590 1959 3620 2011
rect 3996 1959 4026 2011
rect 4198 1959 4228 2011
rect 4636 1959 4666 2011
rect 4838 1959 4868 2011
rect 5244 1959 5274 2011
rect 5446 1959 5476 2011
rect 5884 1959 5914 2011
rect 6086 1959 6116 2011
rect 1615 1604 1667 1610
rect 1615 1546 1667 1552
rect 2205 1604 2257 1610
rect 2205 1546 2257 1552
rect 2863 1604 2915 1610
rect 2863 1546 2915 1552
rect 3453 1604 3505 1610
rect 3453 1546 3505 1552
rect 4111 1604 4163 1610
rect 4111 1546 4163 1552
rect 4701 1604 4753 1610
rect 4701 1546 4753 1552
rect 5359 1604 5411 1610
rect 5359 1546 5411 1552
rect 5949 1604 6001 1610
rect 5949 1546 6001 1552
rect 1604 1167 1656 1173
rect 1604 1109 1656 1115
rect 2216 1167 2268 1173
rect 2216 1109 2268 1115
rect 2852 1167 2904 1173
rect 2852 1109 2904 1115
rect 3464 1167 3516 1173
rect 3464 1109 3516 1115
rect 4100 1167 4152 1173
rect 4100 1109 4152 1115
rect 4712 1167 4764 1173
rect 4712 1109 4764 1115
rect 5348 1167 5400 1173
rect 5348 1109 5400 1115
rect 5960 1167 6012 1173
rect 5960 1109 6012 1115
rect 1725 836 1777 842
rect 1725 778 1777 784
rect 2095 836 2147 842
rect 2095 778 2147 784
rect 2973 836 3025 842
rect 2973 778 3025 784
rect 3343 836 3395 842
rect 3343 778 3395 784
rect 4221 836 4273 842
rect 4221 778 4273 784
rect 4591 836 4643 842
rect 4591 778 4643 784
rect 5469 836 5521 842
rect 5469 778 5521 784
rect 5839 836 5891 842
rect 5839 778 5891 784
rect 1610 633 1662 639
rect 1610 575 1662 581
rect 2210 633 2262 639
rect 2210 575 2262 581
rect 2858 633 2910 639
rect 2858 575 2910 581
rect 3458 633 3510 639
rect 3458 575 3510 581
rect 4106 633 4158 639
rect 4106 575 4158 581
rect 4706 633 4758 639
rect 4706 575 4758 581
rect 5354 633 5406 639
rect 5354 575 5406 581
rect 5954 633 6006 639
rect 5954 575 6006 581
rect 1624 217 1676 223
rect 1624 159 1676 165
rect 2196 217 2248 223
rect 2196 159 2248 165
rect 2872 217 2924 223
rect 2872 159 2924 165
rect 3444 217 3496 223
rect 3444 159 3496 165
rect 4120 217 4172 223
rect 4120 159 4172 165
rect 4692 217 4744 223
rect 4692 159 4744 165
rect 5368 217 5420 223
rect 5368 159 5420 165
rect 5940 217 5992 223
rect 5940 159 5992 165
rect 1473 94 2498 128
rect 2721 94 3746 128
rect 3969 94 4994 128
rect 5217 94 6242 128
rect 1629 4 1689 60
rect 2183 4 2243 60
rect 2877 4 2937 60
rect 3431 4 3491 60
rect 4125 4 4185 60
rect 4679 4 4739 60
rect 5373 4 5433 60
rect 5927 4 5987 60
<< via1 >>
rect 1615 1552 1667 1604
rect 2205 1552 2257 1604
rect 2863 1552 2915 1604
rect 3453 1552 3505 1604
rect 4111 1552 4163 1604
rect 4701 1552 4753 1604
rect 5359 1552 5411 1604
rect 5949 1552 6001 1604
rect 1604 1115 1656 1167
rect 2216 1115 2268 1167
rect 2852 1115 2904 1167
rect 3464 1115 3516 1167
rect 4100 1115 4152 1167
rect 4712 1115 4764 1167
rect 5348 1115 5400 1167
rect 5960 1115 6012 1167
rect 1725 784 1777 836
rect 2095 784 2147 836
rect 2973 784 3025 836
rect 3343 784 3395 836
rect 4221 784 4273 836
rect 4591 784 4643 836
rect 5469 784 5521 836
rect 5839 784 5891 836
rect 1610 581 1662 633
rect 2210 581 2262 633
rect 2858 581 2910 633
rect 3458 581 3510 633
rect 4106 581 4158 633
rect 4706 581 4758 633
rect 5354 581 5406 633
rect 5954 581 6006 633
rect 1624 165 1676 217
rect 2196 165 2248 217
rect 2872 165 2924 217
rect 3444 165 3496 217
rect 4120 165 4172 217
rect 4692 165 4744 217
rect 5368 165 5420 217
rect 5940 165 5992 217
<< metal2 >>
rect 1613 1606 1669 1615
rect 1613 1541 1669 1550
rect 2203 1606 2259 1615
rect 2203 1541 2259 1550
rect 2861 1606 2917 1615
rect 2861 1541 2917 1550
rect 3451 1606 3507 1615
rect 3451 1541 3507 1550
rect 4109 1606 4165 1615
rect 4109 1541 4165 1550
rect 4699 1606 4755 1615
rect 4699 1541 4755 1550
rect 5357 1606 5413 1615
rect 5357 1541 5413 1550
rect 5947 1606 6003 1615
rect 5947 1541 6003 1550
rect 1602 1169 1658 1178
rect 1602 1104 1658 1113
rect 2214 1169 2270 1178
rect 2214 1104 2270 1113
rect 2850 1169 2906 1178
rect 2850 1104 2906 1113
rect 3462 1169 3518 1178
rect 3462 1104 3518 1113
rect 4098 1169 4154 1178
rect 4098 1104 4154 1113
rect 4710 1169 4766 1178
rect 4710 1104 4766 1113
rect 5346 1169 5402 1178
rect 5346 1104 5402 1113
rect 5958 1169 6014 1178
rect 5958 1104 6014 1113
rect 1723 837 1779 846
rect 1723 772 1779 781
rect 2093 837 2149 846
rect 2093 772 2149 781
rect 2971 837 3027 846
rect 2971 772 3027 781
rect 3341 837 3397 846
rect 3341 772 3397 781
rect 4219 837 4275 846
rect 4219 772 4275 781
rect 4589 837 4645 846
rect 4589 772 4645 781
rect 5467 837 5523 846
rect 5467 772 5523 781
rect 5837 837 5893 846
rect 5837 772 5893 781
rect 1608 635 1664 644
rect 1608 570 1664 579
rect 2208 635 2264 644
rect 2208 570 2264 579
rect 2856 635 2912 644
rect 2856 570 2912 579
rect 3456 635 3512 644
rect 3456 570 3512 579
rect 4104 635 4160 644
rect 4104 570 4160 579
rect 4704 635 4760 644
rect 4704 570 4760 579
rect 5352 635 5408 644
rect 5352 570 5408 579
rect 5952 635 6008 644
rect 5952 570 6008 579
rect 1622 219 1678 228
rect 1622 154 1678 163
rect 2194 219 2250 228
rect 2194 154 2250 163
rect 2870 219 2926 228
rect 2870 154 2926 163
rect 3442 219 3498 228
rect 3442 154 3498 163
rect 4118 219 4174 228
rect 4118 154 4174 163
rect 4690 219 4746 228
rect 4690 154 4746 163
rect 5366 219 5422 228
rect 5366 154 5422 163
rect 5938 219 5994 228
rect 5938 154 5994 163
<< via2 >>
rect 1613 1604 1669 1606
rect 1613 1552 1615 1604
rect 1615 1552 1667 1604
rect 1667 1552 1669 1604
rect 1613 1550 1669 1552
rect 2203 1604 2259 1606
rect 2203 1552 2205 1604
rect 2205 1552 2257 1604
rect 2257 1552 2259 1604
rect 2203 1550 2259 1552
rect 2861 1604 2917 1606
rect 2861 1552 2863 1604
rect 2863 1552 2915 1604
rect 2915 1552 2917 1604
rect 2861 1550 2917 1552
rect 3451 1604 3507 1606
rect 3451 1552 3453 1604
rect 3453 1552 3505 1604
rect 3505 1552 3507 1604
rect 3451 1550 3507 1552
rect 4109 1604 4165 1606
rect 4109 1552 4111 1604
rect 4111 1552 4163 1604
rect 4163 1552 4165 1604
rect 4109 1550 4165 1552
rect 4699 1604 4755 1606
rect 4699 1552 4701 1604
rect 4701 1552 4753 1604
rect 4753 1552 4755 1604
rect 4699 1550 4755 1552
rect 5357 1604 5413 1606
rect 5357 1552 5359 1604
rect 5359 1552 5411 1604
rect 5411 1552 5413 1604
rect 5357 1550 5413 1552
rect 5947 1604 6003 1606
rect 5947 1552 5949 1604
rect 5949 1552 6001 1604
rect 6001 1552 6003 1604
rect 5947 1550 6003 1552
rect 1602 1167 1658 1169
rect 1602 1115 1604 1167
rect 1604 1115 1656 1167
rect 1656 1115 1658 1167
rect 1602 1113 1658 1115
rect 2214 1167 2270 1169
rect 2214 1115 2216 1167
rect 2216 1115 2268 1167
rect 2268 1115 2270 1167
rect 2214 1113 2270 1115
rect 2850 1167 2906 1169
rect 2850 1115 2852 1167
rect 2852 1115 2904 1167
rect 2904 1115 2906 1167
rect 2850 1113 2906 1115
rect 3462 1167 3518 1169
rect 3462 1115 3464 1167
rect 3464 1115 3516 1167
rect 3516 1115 3518 1167
rect 3462 1113 3518 1115
rect 4098 1167 4154 1169
rect 4098 1115 4100 1167
rect 4100 1115 4152 1167
rect 4152 1115 4154 1167
rect 4098 1113 4154 1115
rect 4710 1167 4766 1169
rect 4710 1115 4712 1167
rect 4712 1115 4764 1167
rect 4764 1115 4766 1167
rect 4710 1113 4766 1115
rect 5346 1167 5402 1169
rect 5346 1115 5348 1167
rect 5348 1115 5400 1167
rect 5400 1115 5402 1167
rect 5346 1113 5402 1115
rect 5958 1167 6014 1169
rect 5958 1115 5960 1167
rect 5960 1115 6012 1167
rect 6012 1115 6014 1167
rect 5958 1113 6014 1115
rect 1723 836 1779 837
rect 1723 784 1725 836
rect 1725 784 1777 836
rect 1777 784 1779 836
rect 1723 781 1779 784
rect 2093 836 2149 837
rect 2093 784 2095 836
rect 2095 784 2147 836
rect 2147 784 2149 836
rect 2093 781 2149 784
rect 2971 836 3027 837
rect 2971 784 2973 836
rect 2973 784 3025 836
rect 3025 784 3027 836
rect 2971 781 3027 784
rect 3341 836 3397 837
rect 3341 784 3343 836
rect 3343 784 3395 836
rect 3395 784 3397 836
rect 3341 781 3397 784
rect 4219 836 4275 837
rect 4219 784 4221 836
rect 4221 784 4273 836
rect 4273 784 4275 836
rect 4219 781 4275 784
rect 4589 836 4645 837
rect 4589 784 4591 836
rect 4591 784 4643 836
rect 4643 784 4645 836
rect 4589 781 4645 784
rect 5467 836 5523 837
rect 5467 784 5469 836
rect 5469 784 5521 836
rect 5521 784 5523 836
rect 5467 781 5523 784
rect 5837 836 5893 837
rect 5837 784 5839 836
rect 5839 784 5891 836
rect 5891 784 5893 836
rect 5837 781 5893 784
rect 1608 633 1664 635
rect 1608 581 1610 633
rect 1610 581 1662 633
rect 1662 581 1664 633
rect 1608 579 1664 581
rect 2208 633 2264 635
rect 2208 581 2210 633
rect 2210 581 2262 633
rect 2262 581 2264 633
rect 2208 579 2264 581
rect 2856 633 2912 635
rect 2856 581 2858 633
rect 2858 581 2910 633
rect 2910 581 2912 633
rect 2856 579 2912 581
rect 3456 633 3512 635
rect 3456 581 3458 633
rect 3458 581 3510 633
rect 3510 581 3512 633
rect 3456 579 3512 581
rect 4104 633 4160 635
rect 4104 581 4106 633
rect 4106 581 4158 633
rect 4158 581 4160 633
rect 4104 579 4160 581
rect 4704 633 4760 635
rect 4704 581 4706 633
rect 4706 581 4758 633
rect 4758 581 4760 633
rect 4704 579 4760 581
rect 5352 633 5408 635
rect 5352 581 5354 633
rect 5354 581 5406 633
rect 5406 581 5408 633
rect 5352 579 5408 581
rect 5952 633 6008 635
rect 5952 581 5954 633
rect 5954 581 6006 633
rect 6006 581 6008 633
rect 5952 579 6008 581
rect 1622 217 1678 219
rect 1622 165 1624 217
rect 1624 165 1676 217
rect 1676 165 1678 217
rect 1622 163 1678 165
rect 2194 217 2250 219
rect 2194 165 2196 217
rect 2196 165 2248 217
rect 2248 165 2250 217
rect 2194 163 2250 165
rect 2870 217 2926 219
rect 2870 165 2872 217
rect 2872 165 2924 217
rect 2924 165 2926 217
rect 2870 163 2926 165
rect 3442 217 3498 219
rect 3442 165 3444 217
rect 3444 165 3496 217
rect 3496 165 3498 217
rect 3442 163 3498 165
rect 4118 217 4174 219
rect 4118 165 4120 217
rect 4120 165 4172 217
rect 4172 165 4174 217
rect 4118 163 4174 165
rect 4690 217 4746 219
rect 4690 165 4692 217
rect 4692 165 4744 217
rect 4744 165 4746 217
rect 4690 163 4746 165
rect 5366 217 5422 219
rect 5366 165 5368 217
rect 5368 165 5420 217
rect 5420 165 5422 217
rect 5366 163 5422 165
rect 5938 217 5994 219
rect 5938 165 5940 217
rect 5940 165 5992 217
rect 5992 165 5994 217
rect 5938 163 5994 165
<< metal3 >>
rect 1592 1606 1690 1627
rect 1592 1550 1613 1606
rect 1669 1550 1690 1606
rect 1592 1529 1690 1550
rect 2182 1606 2280 1627
rect 2182 1550 2203 1606
rect 2259 1550 2280 1606
rect 2182 1529 2280 1550
rect 2840 1606 2938 1627
rect 2840 1550 2861 1606
rect 2917 1550 2938 1606
rect 2840 1529 2938 1550
rect 3430 1606 3528 1627
rect 3430 1550 3451 1606
rect 3507 1550 3528 1606
rect 3430 1529 3528 1550
rect 4088 1606 4186 1627
rect 4088 1550 4109 1606
rect 4165 1550 4186 1606
rect 4088 1529 4186 1550
rect 4678 1606 4776 1627
rect 4678 1550 4699 1606
rect 4755 1550 4776 1606
rect 4678 1529 4776 1550
rect 5336 1606 5434 1627
rect 5336 1550 5357 1606
rect 5413 1550 5434 1606
rect 5336 1529 5434 1550
rect 5926 1606 6024 1627
rect 5926 1550 5947 1606
rect 6003 1550 6024 1606
rect 5926 1529 6024 1550
rect 1581 1169 1679 1190
rect 1581 1113 1602 1169
rect 1658 1113 1679 1169
rect 1581 1092 1679 1113
rect 2193 1169 2291 1190
rect 2193 1113 2214 1169
rect 2270 1113 2291 1169
rect 2193 1092 2291 1113
rect 2829 1169 2927 1190
rect 2829 1113 2850 1169
rect 2906 1113 2927 1169
rect 2829 1092 2927 1113
rect 3441 1169 3539 1190
rect 3441 1113 3462 1169
rect 3518 1113 3539 1169
rect 3441 1092 3539 1113
rect 4077 1169 4175 1190
rect 4077 1113 4098 1169
rect 4154 1113 4175 1169
rect 4077 1092 4175 1113
rect 4689 1169 4787 1190
rect 4689 1113 4710 1169
rect 4766 1113 4787 1169
rect 4689 1092 4787 1113
rect 5325 1169 5423 1190
rect 5325 1113 5346 1169
rect 5402 1113 5423 1169
rect 5325 1092 5423 1113
rect 5937 1169 6035 1190
rect 5937 1113 5958 1169
rect 6014 1113 6035 1169
rect 5937 1092 6035 1113
rect 1702 837 1800 858
rect 1702 781 1723 837
rect 1779 781 1800 837
rect 1702 760 1800 781
rect 2072 837 2170 858
rect 2072 781 2093 837
rect 2149 781 2170 837
rect 2072 760 2170 781
rect 2950 837 3048 858
rect 2950 781 2971 837
rect 3027 781 3048 837
rect 2950 760 3048 781
rect 3320 837 3418 858
rect 3320 781 3341 837
rect 3397 781 3418 837
rect 3320 760 3418 781
rect 4198 837 4296 858
rect 4198 781 4219 837
rect 4275 781 4296 837
rect 4198 760 4296 781
rect 4568 837 4666 858
rect 4568 781 4589 837
rect 4645 781 4666 837
rect 4568 760 4666 781
rect 5446 837 5544 858
rect 5446 781 5467 837
rect 5523 781 5544 837
rect 5446 760 5544 781
rect 5816 837 5914 858
rect 5816 781 5837 837
rect 5893 781 5914 837
rect 5816 760 5914 781
rect 1587 635 1685 656
rect 1587 579 1608 635
rect 1664 579 1685 635
rect 1587 558 1685 579
rect 2187 635 2285 656
rect 2187 579 2208 635
rect 2264 579 2285 635
rect 2187 558 2285 579
rect 2835 635 2933 656
rect 2835 579 2856 635
rect 2912 579 2933 635
rect 2835 558 2933 579
rect 3435 635 3533 656
rect 3435 579 3456 635
rect 3512 579 3533 635
rect 3435 558 3533 579
rect 4083 635 4181 656
rect 4083 579 4104 635
rect 4160 579 4181 635
rect 4083 558 4181 579
rect 4683 635 4781 656
rect 4683 579 4704 635
rect 4760 579 4781 635
rect 4683 558 4781 579
rect 5331 635 5429 656
rect 5331 579 5352 635
rect 5408 579 5429 635
rect 5331 558 5429 579
rect 5931 635 6029 656
rect 5931 579 5952 635
rect 6008 579 6029 635
rect 5931 558 6029 579
rect 1601 219 1699 240
rect 1601 163 1622 219
rect 1678 163 1699 219
rect 1601 142 1699 163
rect 2173 219 2271 240
rect 2173 163 2194 219
rect 2250 163 2271 219
rect 2173 142 2271 163
rect 2849 219 2947 240
rect 2849 163 2870 219
rect 2926 163 2947 219
rect 2849 142 2947 163
rect 3421 219 3519 240
rect 3421 163 3442 219
rect 3498 163 3519 219
rect 3421 142 3519 163
rect 4097 219 4195 240
rect 4097 163 4118 219
rect 4174 163 4195 219
rect 4097 142 4195 163
rect 4669 219 4767 240
rect 4669 163 4690 219
rect 4746 163 4767 219
rect 4669 142 4767 163
rect 5345 219 5443 240
rect 5345 163 5366 219
rect 5422 163 5443 219
rect 5345 142 5443 163
rect 5917 219 6015 240
rect 5917 163 5938 219
rect 5994 163 6015 219
rect 5917 142 6015 163
use contact_23  contact_23_0
timestamp 1634918361
transform 1 0 5942 0 1 1541
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1634918361
transform 1 0 5949 0 1 1546
box 0 0 1 1
use contact_23  contact_23_1
timestamp 1634918361
transform 1 0 5832 0 1 772
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1634918361
transform 1 0 5839 0 1 778
box 0 0 1 1
use contact_23  contact_23_2
timestamp 1634918361
transform 1 0 5947 0 1 570
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1634918361
transform 1 0 5954 0 1 575
box 0 0 1 1
use contact_23  contact_23_3
timestamp 1634918361
transform 1 0 5953 0 1 1104
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1634918361
transform 1 0 5960 0 1 1109
box 0 0 1 1
use contact_23  contact_23_4
timestamp 1634918361
transform 1 0 5933 0 1 154
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1634918361
transform 1 0 5940 0 1 159
box 0 0 1 1
use contact_23  contact_23_5
timestamp 1634918361
transform 1 0 5352 0 1 1541
box 0 0 1 1
use contact_22  contact_22_5
timestamp 1634918361
transform 1 0 5359 0 1 1546
box 0 0 1 1
use contact_23  contact_23_6
timestamp 1634918361
transform 1 0 5462 0 1 772
box 0 0 1 1
use contact_22  contact_22_6
timestamp 1634918361
transform 1 0 5469 0 1 778
box 0 0 1 1
use contact_23  contact_23_7
timestamp 1634918361
transform 1 0 5347 0 1 570
box 0 0 1 1
use contact_22  contact_22_7
timestamp 1634918361
transform 1 0 5354 0 1 575
box 0 0 1 1
use contact_23  contact_23_8
timestamp 1634918361
transform 1 0 5341 0 1 1104
box 0 0 1 1
use contact_22  contact_22_8
timestamp 1634918361
transform 1 0 5348 0 1 1109
box 0 0 1 1
use contact_23  contact_23_9
timestamp 1634918361
transform 1 0 5361 0 1 154
box 0 0 1 1
use contact_22  contact_22_9
timestamp 1634918361
transform 1 0 5368 0 1 159
box 0 0 1 1
use contact_23  contact_23_10
timestamp 1634918361
transform 1 0 4694 0 1 1541
box 0 0 1 1
use contact_22  contact_22_10
timestamp 1634918361
transform 1 0 4701 0 1 1546
box 0 0 1 1
use contact_23  contact_23_11
timestamp 1634918361
transform 1 0 4584 0 1 772
box 0 0 1 1
use contact_22  contact_22_11
timestamp 1634918361
transform 1 0 4591 0 1 778
box 0 0 1 1
use contact_23  contact_23_12
timestamp 1634918361
transform 1 0 4699 0 1 570
box 0 0 1 1
use contact_22  contact_22_12
timestamp 1634918361
transform 1 0 4706 0 1 575
box 0 0 1 1
use contact_23  contact_23_13
timestamp 1634918361
transform 1 0 4705 0 1 1104
box 0 0 1 1
use contact_22  contact_22_13
timestamp 1634918361
transform 1 0 4712 0 1 1109
box 0 0 1 1
use contact_23  contact_23_14
timestamp 1634918361
transform 1 0 4685 0 1 154
box 0 0 1 1
use contact_22  contact_22_14
timestamp 1634918361
transform 1 0 4692 0 1 159
box 0 0 1 1
use contact_23  contact_23_15
timestamp 1634918361
transform 1 0 4104 0 1 1541
box 0 0 1 1
use contact_22  contact_22_15
timestamp 1634918361
transform 1 0 4111 0 1 1546
box 0 0 1 1
use contact_23  contact_23_16
timestamp 1634918361
transform 1 0 4214 0 1 772
box 0 0 1 1
use contact_22  contact_22_16
timestamp 1634918361
transform 1 0 4221 0 1 778
box 0 0 1 1
use contact_23  contact_23_17
timestamp 1634918361
transform 1 0 4099 0 1 570
box 0 0 1 1
use contact_22  contact_22_17
timestamp 1634918361
transform 1 0 4106 0 1 575
box 0 0 1 1
use contact_23  contact_23_18
timestamp 1634918361
transform 1 0 4093 0 1 1104
box 0 0 1 1
use contact_22  contact_22_18
timestamp 1634918361
transform 1 0 4100 0 1 1109
box 0 0 1 1
use contact_23  contact_23_19
timestamp 1634918361
transform 1 0 4113 0 1 154
box 0 0 1 1
use contact_22  contact_22_19
timestamp 1634918361
transform 1 0 4120 0 1 159
box 0 0 1 1
use contact_23  contact_23_20
timestamp 1634918361
transform 1 0 3446 0 1 1541
box 0 0 1 1
use contact_22  contact_22_20
timestamp 1634918361
transform 1 0 3453 0 1 1546
box 0 0 1 1
use contact_23  contact_23_21
timestamp 1634918361
transform 1 0 3336 0 1 772
box 0 0 1 1
use contact_22  contact_22_21
timestamp 1634918361
transform 1 0 3343 0 1 778
box 0 0 1 1
use contact_23  contact_23_22
timestamp 1634918361
transform 1 0 3451 0 1 570
box 0 0 1 1
use contact_22  contact_22_22
timestamp 1634918361
transform 1 0 3458 0 1 575
box 0 0 1 1
use contact_23  contact_23_23
timestamp 1634918361
transform 1 0 3457 0 1 1104
box 0 0 1 1
use contact_22  contact_22_23
timestamp 1634918361
transform 1 0 3464 0 1 1109
box 0 0 1 1
use contact_23  contact_23_24
timestamp 1634918361
transform 1 0 3437 0 1 154
box 0 0 1 1
use contact_22  contact_22_24
timestamp 1634918361
transform 1 0 3444 0 1 159
box 0 0 1 1
use contact_23  contact_23_25
timestamp 1634918361
transform 1 0 2856 0 1 1541
box 0 0 1 1
use contact_22  contact_22_25
timestamp 1634918361
transform 1 0 2863 0 1 1546
box 0 0 1 1
use contact_23  contact_23_26
timestamp 1634918361
transform 1 0 2966 0 1 772
box 0 0 1 1
use contact_22  contact_22_26
timestamp 1634918361
transform 1 0 2973 0 1 778
box 0 0 1 1
use contact_23  contact_23_27
timestamp 1634918361
transform 1 0 2851 0 1 570
box 0 0 1 1
use contact_22  contact_22_27
timestamp 1634918361
transform 1 0 2858 0 1 575
box 0 0 1 1
use contact_23  contact_23_28
timestamp 1634918361
transform 1 0 2845 0 1 1104
box 0 0 1 1
use contact_22  contact_22_28
timestamp 1634918361
transform 1 0 2852 0 1 1109
box 0 0 1 1
use contact_23  contact_23_29
timestamp 1634918361
transform 1 0 2865 0 1 154
box 0 0 1 1
use contact_22  contact_22_29
timestamp 1634918361
transform 1 0 2872 0 1 159
box 0 0 1 1
use contact_23  contact_23_30
timestamp 1634918361
transform 1 0 2198 0 1 1541
box 0 0 1 1
use contact_22  contact_22_30
timestamp 1634918361
transform 1 0 2205 0 1 1546
box 0 0 1 1
use contact_23  contact_23_31
timestamp 1634918361
transform 1 0 2088 0 1 772
box 0 0 1 1
use contact_22  contact_22_31
timestamp 1634918361
transform 1 0 2095 0 1 778
box 0 0 1 1
use contact_23  contact_23_32
timestamp 1634918361
transform 1 0 2203 0 1 570
box 0 0 1 1
use contact_22  contact_22_32
timestamp 1634918361
transform 1 0 2210 0 1 575
box 0 0 1 1
use contact_23  contact_23_33
timestamp 1634918361
transform 1 0 2209 0 1 1104
box 0 0 1 1
use contact_22  contact_22_33
timestamp 1634918361
transform 1 0 2216 0 1 1109
box 0 0 1 1
use contact_23  contact_23_34
timestamp 1634918361
transform 1 0 2189 0 1 154
box 0 0 1 1
use contact_22  contact_22_34
timestamp 1634918361
transform 1 0 2196 0 1 159
box 0 0 1 1
use contact_23  contact_23_35
timestamp 1634918361
transform 1 0 1608 0 1 1541
box 0 0 1 1
use contact_22  contact_22_35
timestamp 1634918361
transform 1 0 1615 0 1 1546
box 0 0 1 1
use contact_23  contact_23_36
timestamp 1634918361
transform 1 0 1718 0 1 772
box 0 0 1 1
use contact_22  contact_22_36
timestamp 1634918361
transform 1 0 1725 0 1 778
box 0 0 1 1
use contact_23  contact_23_37
timestamp 1634918361
transform 1 0 1603 0 1 570
box 0 0 1 1
use contact_22  contact_22_37
timestamp 1634918361
transform 1 0 1610 0 1 575
box 0 0 1 1
use contact_23  contact_23_38
timestamp 1634918361
transform 1 0 1597 0 1 1104
box 0 0 1 1
use contact_22  contact_22_38
timestamp 1634918361
transform 1 0 1604 0 1 1109
box 0 0 1 1
use contact_23  contact_23_39
timestamp 1634918361
transform 1 0 1617 0 1 154
box 0 0 1 1
use contact_22  contact_22_39
timestamp 1634918361
transform 1 0 1624 0 1 159
box 0 0 1 1
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_0
timestamp 1634918361
transform -1 0 6242 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_1
timestamp 1634918361
transform 1 0 5118 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_2
timestamp 1634918361
transform -1 0 4994 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_3
timestamp 1634918361
transform 1 0 3870 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_4
timestamp 1634918361
transform -1 0 3746 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_5
timestamp 1634918361
transform 1 0 2622 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_6
timestamp 1634918361
transform -1 0 2498 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_7
timestamp 1634918361
transform 1 0 1374 0 1 0
box -376 4 880 2011
<< labels >>
rlabel metal1 s 1629 4 1689 60 4 data_0
port 1 nsew
rlabel metal1 s 1500 1959 1530 2011 4 bl_0
port 2 nsew
rlabel metal1 s 1702 1959 1732 2011 4 br_0
port 3 nsew
rlabel metal3 s 2849 142 2947 240 4 vdd
port 4 nsew
rlabel metal3 s 2193 1092 2291 1190 4 vdd
port 4 nsew
rlabel metal3 s 2829 1092 2927 1190 4 vdd
port 4 nsew
rlabel metal3 s 3421 142 3519 240 4 vdd
port 4 nsew
rlabel metal3 s 4689 1092 4787 1190 4 vdd
port 4 nsew
rlabel metal3 s 1601 142 1699 240 4 vdd
port 4 nsew
rlabel metal3 s 4077 1092 4175 1190 4 vdd
port 4 nsew
rlabel metal3 s 5345 142 5443 240 4 vdd
port 4 nsew
rlabel metal3 s 5325 1092 5423 1190 4 vdd
port 4 nsew
rlabel metal3 s 4669 142 4767 240 4 vdd
port 4 nsew
rlabel metal3 s 3441 1092 3539 1190 4 vdd
port 4 nsew
rlabel metal3 s 2173 142 2271 240 4 vdd
port 4 nsew
rlabel metal3 s 4097 142 4195 240 4 vdd
port 4 nsew
rlabel metal3 s 1581 1092 1679 1190 4 vdd
port 4 nsew
rlabel metal3 s 5917 142 6015 240 4 vdd
port 4 nsew
rlabel metal3 s 5937 1092 6035 1190 4 vdd
port 4 nsew
rlabel metal3 s 2187 558 2285 656 4 gnd
port 5 nsew
rlabel metal3 s 5336 1529 5434 1627 4 gnd
port 5 nsew
rlabel metal3 s 2072 760 2170 858 4 gnd
port 5 nsew
rlabel metal3 s 3320 760 3418 858 4 gnd
port 5 nsew
rlabel metal3 s 1592 1529 1690 1627 4 gnd
port 5 nsew
rlabel metal3 s 2950 760 3048 858 4 gnd
port 5 nsew
rlabel metal3 s 5331 558 5429 656 4 gnd
port 5 nsew
rlabel metal3 s 3430 1529 3528 1627 4 gnd
port 5 nsew
rlabel metal3 s 4678 1529 4776 1627 4 gnd
port 5 nsew
rlabel metal3 s 5816 760 5914 858 4 gnd
port 5 nsew
rlabel metal3 s 4568 760 4666 858 4 gnd
port 5 nsew
rlabel metal3 s 1587 558 1685 656 4 gnd
port 5 nsew
rlabel metal3 s 1702 760 1800 858 4 gnd
port 5 nsew
rlabel metal3 s 5931 558 6029 656 4 gnd
port 5 nsew
rlabel metal3 s 4083 558 4181 656 4 gnd
port 5 nsew
rlabel metal3 s 4088 1529 4186 1627 4 gnd
port 5 nsew
rlabel metal3 s 3435 558 3533 656 4 gnd
port 5 nsew
rlabel metal3 s 2182 1529 2280 1627 4 gnd
port 5 nsew
rlabel metal3 s 4198 760 4296 858 4 gnd
port 5 nsew
rlabel metal3 s 5446 760 5544 858 4 gnd
port 5 nsew
rlabel metal3 s 5926 1529 6024 1627 4 gnd
port 5 nsew
rlabel metal3 s 4683 558 4781 656 4 gnd
port 5 nsew
rlabel metal3 s 2840 1529 2938 1627 4 gnd
port 5 nsew
rlabel metal3 s 2835 558 2933 656 4 gnd
port 5 nsew
rlabel metal1 s 2183 4 2243 60 4 data_1
port 6 nsew
rlabel metal1 s 2342 1959 2372 2011 4 bl_1
port 7 nsew
rlabel metal1 s 2140 1959 2170 2011 4 br_1
port 8 nsew
rlabel metal1 s 2877 4 2937 60 4 data_2
port 9 nsew
rlabel metal1 s 2748 1959 2778 2011 4 bl_2
port 10 nsew
rlabel metal1 s 2950 1959 2980 2011 4 br_2
port 11 nsew
rlabel metal1 s 3431 4 3491 60 4 data_3
port 12 nsew
rlabel metal1 s 3590 1959 3620 2011 4 bl_3
port 13 nsew
rlabel metal1 s 3388 1959 3418 2011 4 br_3
port 14 nsew
rlabel metal1 s 4125 4 4185 60 4 data_4
port 15 nsew
rlabel metal1 s 3996 1959 4026 2011 4 bl_4
port 16 nsew
rlabel metal1 s 4198 1959 4228 2011 4 br_4
port 17 nsew
rlabel metal1 s 4679 4 4739 60 4 data_5
port 18 nsew
rlabel metal1 s 4838 1959 4868 2011 4 bl_5
port 19 nsew
rlabel metal1 s 4636 1959 4666 2011 4 br_5
port 20 nsew
rlabel metal1 s 5373 4 5433 60 4 data_6
port 21 nsew
rlabel metal1 s 5244 1959 5274 2011 4 bl_6
port 22 nsew
rlabel metal1 s 5446 1959 5476 2011 4 br_6
port 23 nsew
rlabel metal1 s 5927 4 5987 60 4 data_7
port 24 nsew
rlabel metal1 s 6086 1959 6116 2011 4 bl_7
port 25 nsew
rlabel metal1 s 5884 1959 5914 2011 4 br_7
port 26 nsew
rlabel metal1 s 1473 94 2498 128 4 en_0
port 27 nsew
rlabel metal1 s 2721 94 3746 128 4 en_1
port 28 nsew
rlabel metal1 s 3969 94 4994 128 4 en_2
port 29 nsew
rlabel metal1 s 5217 94 6242 128 4 en_3
port 30 nsew
<< properties >>
string FIXED_BBOX 0 0 6242 2011
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 855314
string GDS_START 836966
<< end >>
