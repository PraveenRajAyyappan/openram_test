magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1235 -1186 1385 1335
<< labels >>
rlabel poly s 75 74 75 74 4 G
port 1 nsew
rlabel mvpsubdiff s 25 74 25 74 4 S
rlabel mvpsubdiff s 125 74 125 74 4 D
<< properties >>
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1131570
string GDS_START 1130922
<< end >>
