magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1296 -1277 4604 2731
<< nwell >>
rect -36 679 3344 1471
<< locali >>
rect 0 1397 3308 1431
rect 64 636 98 702
rect 179 653 449 687
rect 551 674 925 708
rect 1241 690 1725 724
rect 2473 690 2507 724
rect 551 670 585 674
rect 0 -17 3308 17
use pinv_12  pinv_12_0
timestamp 1634918361
transform 1 0 1644 0 1 0
box -36 -17 1700 1471
use pinv_6  pinv_6_0
timestamp 1634918361
transform 1 0 844 0 1 0
box -36 -17 836 1471
use pinv_5  pinv_5_0
timestamp 1634918361
transform 1 0 368 0 1 0
box -36 -17 512 1471
use pinv_4  pinv_4_0
timestamp 1634918361
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 2490 707 2490 707 4 Z
port 1 nsew
rlabel locali s 81 669 81 669 4 A
port 2 nsew
rlabel locali s 1654 0 1654 0 4 gnd
port 3 nsew
rlabel locali s 1654 1414 1654 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 3308 1414
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1198328
string GDS_START 1196846
<< end >>
