magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1260 -1316 7143 7636
<< locali >>
rect 5288 6183 5865 6217
rect 4148 6112 4164 6146
rect 4198 6112 4367 6146
rect 3828 6004 3844 6038
rect 3878 6004 4367 6038
rect 3748 5812 3764 5846
rect 3798 5812 4367 5846
rect 4148 5704 4164 5738
rect 4198 5704 4367 5738
rect 5288 5633 5865 5667
rect 5288 5393 5865 5427
rect 4148 5322 4164 5356
rect 4198 5322 4367 5356
rect 3668 5214 3684 5248
rect 3718 5214 4367 5248
rect 3588 5022 3604 5056
rect 3638 5022 4367 5056
rect 4148 4914 4164 4948
rect 4198 4914 4367 4948
rect 5288 4843 5865 4877
rect 5288 4603 5865 4637
rect 4068 4532 4084 4566
rect 4118 4532 4367 4566
rect 3828 4424 3844 4458
rect 3878 4424 4367 4458
rect 3748 4232 3764 4266
rect 3798 4232 4367 4266
rect 4068 4124 4084 4158
rect 4118 4124 4367 4158
rect 5288 4053 5865 4087
rect 3510 3847 3544 3863
rect 5288 3813 5865 3847
rect 3510 3797 3544 3813
rect 4068 3742 4084 3776
rect 4118 3742 4367 3776
rect 3668 3634 3684 3668
rect 3718 3634 4367 3668
rect 3588 3442 3604 3476
rect 3638 3442 4367 3476
rect 4068 3334 4084 3368
rect 4118 3334 4367 3368
rect 3510 3297 3544 3313
rect 5288 3263 5865 3297
rect 3510 3247 3544 3263
rect 3510 3057 3544 3073
rect 5288 3023 5865 3057
rect 524 3007 558 3023
rect 3510 3007 3544 3023
rect 240 2973 256 3007
rect 290 2973 524 3007
rect 524 2957 558 2973
rect 3988 2952 4004 2986
rect 4038 2952 4367 2986
rect 3828 2844 3844 2878
rect 3878 2844 4367 2878
rect 3748 2652 3764 2686
rect 3798 2652 4367 2686
rect 444 2557 478 2573
rect 160 2523 176 2557
rect 210 2523 444 2557
rect 3988 2544 4004 2578
rect 4038 2544 4367 2578
rect 444 2507 478 2523
rect 3510 2507 3544 2523
rect 5288 2473 5865 2507
rect 3510 2457 3544 2473
rect 5288 2233 5865 2267
rect 3988 2162 4004 2196
rect 4038 2162 4367 2196
rect 3668 2054 3684 2088
rect 3718 2054 4367 2088
rect 3588 1862 3604 1896
rect 3638 1862 4367 1896
rect 3988 1754 4004 1788
rect 4038 1754 4367 1788
rect 5288 1683 5865 1717
rect 3510 1477 3544 1493
rect 5288 1443 5865 1477
rect 3510 1427 3544 1443
rect 3908 1372 3924 1406
rect 3958 1372 4367 1406
rect 3828 1264 3844 1298
rect 3878 1264 4367 1298
rect 3748 1072 3764 1106
rect 3798 1072 4367 1106
rect 3908 964 3924 998
rect 3958 964 4367 998
rect 3510 927 3544 943
rect 5288 893 5865 927
rect 3510 877 3544 893
rect 3510 687 3544 703
rect 5288 653 5865 687
rect 524 637 558 653
rect 3510 637 3544 653
rect 80 603 96 637
rect 130 603 524 637
rect 524 587 558 603
rect 3908 582 3924 616
rect 3958 582 4367 616
rect 3668 474 3684 508
rect 3718 474 4367 508
rect 3588 282 3604 316
rect 3638 282 4367 316
rect 444 187 478 203
rect 0 153 16 187
rect 50 153 444 187
rect 3908 174 3924 208
rect 3958 174 4367 208
rect 444 137 478 153
rect 3510 137 3544 153
rect 5288 103 5865 137
rect 3510 87 3544 103
<< viali >>
rect 4164 6112 4198 6146
rect 3844 6004 3878 6038
rect 3764 5812 3798 5846
rect 4164 5704 4198 5738
rect 4164 5322 4198 5356
rect 3684 5214 3718 5248
rect 3604 5022 3638 5056
rect 4164 4914 4198 4948
rect 4084 4532 4118 4566
rect 3844 4424 3878 4458
rect 3764 4232 3798 4266
rect 4084 4124 4118 4158
rect 3510 3813 3544 3847
rect 4084 3742 4118 3776
rect 3684 3634 3718 3668
rect 3604 3442 3638 3476
rect 4084 3334 4118 3368
rect 3510 3263 3544 3297
rect 3510 3023 3544 3057
rect 256 2973 290 3007
rect 524 2973 558 3007
rect 4004 2952 4038 2986
rect 3844 2844 3878 2878
rect 3764 2652 3798 2686
rect 176 2523 210 2557
rect 444 2523 478 2557
rect 4004 2544 4038 2578
rect 3510 2473 3544 2507
rect 4004 2162 4038 2196
rect 3684 2054 3718 2088
rect 3604 1862 3638 1896
rect 4004 1754 4038 1788
rect 3510 1443 3544 1477
rect 3924 1372 3958 1406
rect 3844 1264 3878 1298
rect 3764 1072 3798 1106
rect 3924 964 3958 998
rect 3510 893 3544 927
rect 3510 653 3544 687
rect 96 603 130 637
rect 524 603 558 637
rect 3924 582 3958 616
rect 3684 474 3718 508
rect 3604 282 3638 316
rect 16 153 50 187
rect 444 153 478 187
rect 3924 174 3958 208
rect 3510 103 3544 137
<< metal1 >>
rect 3607 5068 3635 6348
rect 3687 5260 3715 6348
rect 3767 5858 3795 6348
rect 3847 6050 3875 6348
rect 3838 6038 3884 6050
rect 3838 6004 3844 6038
rect 3878 6004 3884 6038
rect 3838 5992 3884 6004
rect 3758 5846 3804 5858
rect 3758 5812 3764 5846
rect 3798 5812 3804 5846
rect 3758 5800 3804 5812
rect 3678 5248 3724 5260
rect 3678 5214 3684 5248
rect 3718 5214 3724 5248
rect 3678 5202 3724 5214
rect 3598 5056 3644 5068
rect 3598 5022 3604 5056
rect 3638 5022 3644 5056
rect 3598 5010 3644 5022
rect 19 199 47 3950
rect 99 649 127 3950
rect 179 2569 207 3950
rect 259 3019 287 3950
rect 3495 3804 3501 3856
rect 3553 3804 3559 3856
rect 3607 3488 3635 5010
rect 3687 3680 3715 5202
rect 3767 4278 3795 5800
rect 3847 4470 3875 5992
rect 3838 4458 3884 4470
rect 3838 4424 3844 4458
rect 3878 4424 3884 4458
rect 3838 4412 3884 4424
rect 3758 4266 3804 4278
rect 3758 4232 3764 4266
rect 3798 4232 3804 4266
rect 3758 4220 3804 4232
rect 3678 3668 3724 3680
rect 3678 3634 3684 3668
rect 3718 3634 3724 3668
rect 3678 3622 3724 3634
rect 3598 3476 3644 3488
rect 3598 3442 3604 3476
rect 3638 3442 3644 3476
rect 3598 3430 3644 3442
rect 3495 3254 3501 3306
rect 3553 3254 3559 3306
rect 250 3007 296 3019
rect 3495 3014 3501 3066
rect 3553 3014 3559 3066
rect 250 2973 256 3007
rect 290 2973 296 3007
rect 250 2961 296 2973
rect 512 3007 570 3013
rect 512 2973 524 3007
rect 558 2973 570 3007
rect 512 2967 570 2973
rect 170 2557 216 2569
rect 170 2523 176 2557
rect 210 2523 216 2557
rect 170 2511 216 2523
rect 90 637 136 649
rect 90 603 96 637
rect 130 603 136 637
rect 90 591 136 603
rect 10 187 56 199
rect 10 153 16 187
rect 50 153 56 187
rect 10 141 56 153
rect 19 0 47 141
rect 99 0 127 591
rect 179 0 207 2511
rect 259 0 287 2961
rect 432 2557 490 2563
rect 432 2523 444 2557
rect 478 2523 490 2557
rect 432 2517 490 2523
rect 3495 2464 3501 2516
rect 3553 2464 3559 2516
rect 3607 1908 3635 3430
rect 3687 2100 3715 3622
rect 3767 2698 3795 4220
rect 3847 2890 3875 4412
rect 3838 2878 3884 2890
rect 3838 2844 3844 2878
rect 3878 2844 3884 2878
rect 3838 2832 3884 2844
rect 3758 2686 3804 2698
rect 3758 2652 3764 2686
rect 3798 2652 3804 2686
rect 3758 2640 3804 2652
rect 3678 2088 3724 2100
rect 3678 2054 3684 2088
rect 3718 2054 3724 2088
rect 3678 2042 3724 2054
rect 3598 1896 3644 1908
rect 3598 1862 3604 1896
rect 3638 1862 3644 1896
rect 3598 1850 3644 1862
rect 3495 1434 3501 1486
rect 3553 1434 3559 1486
rect 3495 884 3501 936
rect 3553 884 3559 936
rect 3495 644 3501 696
rect 3553 644 3559 696
rect 512 637 570 643
rect 512 603 524 637
rect 558 603 570 637
rect 512 597 570 603
rect 3607 328 3635 1850
rect 3687 520 3715 2042
rect 3767 1118 3795 2640
rect 3847 1310 3875 2832
rect 3927 2402 3955 6348
rect 4007 2998 4035 6348
rect 4087 4578 4115 6348
rect 4167 6158 4195 6348
rect 4158 6146 4204 6158
rect 4158 6112 4164 6146
rect 4198 6112 4204 6146
rect 4158 6100 4204 6112
rect 4167 5750 4195 6100
rect 4493 5958 4541 6290
rect 4917 5958 4967 6288
rect 4485 5906 4491 5958
rect 4543 5906 4549 5958
rect 4910 5906 4916 5958
rect 4968 5906 4974 5958
rect 5307 5951 5335 6320
rect 5703 5951 5731 6320
rect 4158 5738 4204 5750
rect 4158 5704 4164 5738
rect 4198 5704 4204 5738
rect 4158 5692 4204 5704
rect 4167 5368 4195 5692
rect 4493 5586 4541 5906
rect 4917 5588 4967 5906
rect 5289 5899 5295 5951
rect 5347 5899 5353 5951
rect 5685 5899 5691 5951
rect 5743 5899 5749 5951
rect 4485 5534 4491 5586
rect 4543 5534 4549 5586
rect 4910 5536 4916 5588
rect 4968 5536 4974 5588
rect 5307 5556 5335 5899
rect 5703 5556 5731 5899
rect 4158 5356 4204 5368
rect 4158 5322 4164 5356
rect 4198 5322 4204 5356
rect 4158 5310 4204 5322
rect 4167 4960 4195 5310
rect 4493 5168 4541 5534
rect 4917 5168 4967 5536
rect 5289 5504 5295 5556
rect 5347 5504 5353 5556
rect 5685 5504 5691 5556
rect 5743 5504 5749 5556
rect 4485 5116 4491 5168
rect 4543 5116 4549 5168
rect 4910 5116 4916 5168
rect 4968 5116 4974 5168
rect 5307 5161 5335 5504
rect 5703 5161 5731 5504
rect 4158 4948 4204 4960
rect 4158 4914 4164 4948
rect 4198 4914 4204 4948
rect 4158 4902 4204 4914
rect 4078 4566 4124 4578
rect 4078 4532 4084 4566
rect 4118 4532 4124 4566
rect 4078 4520 4124 4532
rect 4087 4170 4115 4520
rect 4078 4158 4124 4170
rect 4078 4124 4084 4158
rect 4118 4124 4124 4158
rect 4078 4112 4124 4124
rect 4087 3788 4115 4112
rect 4078 3776 4124 3788
rect 4078 3742 4084 3776
rect 4118 3742 4124 3776
rect 4078 3730 4124 3742
rect 4087 3380 4115 3730
rect 4167 3587 4195 4902
rect 4493 4796 4541 5116
rect 4917 4798 4967 5116
rect 5289 5109 5295 5161
rect 5347 5109 5353 5161
rect 5685 5109 5691 5161
rect 5743 5109 5749 5161
rect 4485 4744 4491 4796
rect 4543 4744 4549 4796
rect 4910 4746 4916 4798
rect 4968 4746 4974 4798
rect 5307 4766 5335 5109
rect 5703 4766 5731 5109
rect 4493 4378 4541 4744
rect 4917 4378 4967 4746
rect 5289 4714 5295 4766
rect 5347 4714 5353 4766
rect 5685 4714 5691 4766
rect 5743 4714 5749 4766
rect 4485 4326 4491 4378
rect 4543 4326 4549 4378
rect 4910 4326 4916 4378
rect 4968 4326 4974 4378
rect 5307 4371 5335 4714
rect 5703 4371 5731 4714
rect 4493 4006 4541 4326
rect 4917 4008 4967 4326
rect 5289 4319 5295 4371
rect 5347 4319 5353 4371
rect 5685 4319 5691 4371
rect 5743 4319 5749 4371
rect 4485 3954 4491 4006
rect 4543 3954 4549 4006
rect 4910 3956 4916 4008
rect 4968 3956 4974 4008
rect 5307 3976 5335 4319
rect 5703 3976 5731 4319
rect 4493 3588 4541 3954
rect 4917 3588 4967 3956
rect 5289 3924 5295 3976
rect 5347 3924 5353 3976
rect 5685 3924 5691 3976
rect 5743 3924 5749 3976
rect 4155 3581 4207 3587
rect 4485 3536 4491 3588
rect 4543 3536 4549 3588
rect 4910 3536 4916 3588
rect 4968 3536 4974 3588
rect 5307 3581 5335 3924
rect 5703 3581 5731 3924
rect 4155 3523 4207 3529
rect 4078 3368 4124 3380
rect 4078 3334 4084 3368
rect 4118 3334 4124 3368
rect 4078 3322 4124 3334
rect 4087 3192 4115 3322
rect 4075 3186 4127 3192
rect 4075 3128 4127 3134
rect 3998 2986 4044 2998
rect 3998 2952 4004 2986
rect 4038 2952 4044 2986
rect 3998 2940 4044 2952
rect 4007 2797 4035 2940
rect 3995 2791 4047 2797
rect 3995 2733 4047 2739
rect 4007 2590 4035 2733
rect 3998 2578 4044 2590
rect 3998 2544 4004 2578
rect 4038 2544 4044 2578
rect 3998 2532 4044 2544
rect 3915 2396 3967 2402
rect 3915 2338 3967 2344
rect 3927 1418 3955 2338
rect 4007 2208 4035 2532
rect 3998 2196 4044 2208
rect 3998 2162 4004 2196
rect 4038 2162 4044 2196
rect 3998 2150 4044 2162
rect 4007 1800 4035 2150
rect 3998 1788 4044 1800
rect 3998 1754 4004 1788
rect 4038 1754 4044 1788
rect 3998 1742 4044 1754
rect 3918 1406 3964 1418
rect 3918 1372 3924 1406
rect 3958 1372 3964 1406
rect 3918 1360 3964 1372
rect 3838 1298 3884 1310
rect 3838 1264 3844 1298
rect 3878 1264 3884 1298
rect 3838 1252 3884 1264
rect 3847 1217 3875 1252
rect 3835 1211 3887 1217
rect 3835 1153 3887 1159
rect 3758 1106 3804 1118
rect 3758 1072 3764 1106
rect 3798 1072 3804 1106
rect 3758 1060 3804 1072
rect 3767 822 3795 1060
rect 3755 816 3807 822
rect 3755 758 3807 764
rect 3678 508 3724 520
rect 3678 474 3684 508
rect 3718 474 3724 508
rect 3678 462 3724 474
rect 3687 427 3715 462
rect 3675 421 3727 427
rect 3675 363 3727 369
rect 3598 316 3644 328
rect 3598 282 3604 316
rect 3638 282 3644 316
rect 3598 270 3644 282
rect 432 187 490 193
rect 432 153 444 187
rect 478 153 490 187
rect 432 147 490 153
rect 3495 94 3501 146
rect 3553 94 3559 146
rect 3607 32 3635 270
rect 3595 26 3647 32
rect 3687 0 3715 363
rect 3767 0 3795 758
rect 3847 0 3875 1153
rect 3927 1010 3955 1360
rect 3918 998 3964 1010
rect 3918 964 3924 998
rect 3958 964 3964 998
rect 3918 952 3964 964
rect 3927 628 3955 952
rect 3918 616 3964 628
rect 3918 582 3924 616
rect 3958 582 3964 616
rect 3918 570 3964 582
rect 3927 220 3955 570
rect 3918 208 3964 220
rect 3918 174 3924 208
rect 3958 174 3964 208
rect 3918 162 3964 174
rect 3927 0 3955 162
rect 4007 0 4035 1742
rect 4087 0 4115 3128
rect 4167 0 4195 3523
rect 4493 3216 4541 3536
rect 4917 3218 4967 3536
rect 5289 3529 5295 3581
rect 5347 3529 5353 3581
rect 5685 3529 5691 3581
rect 5743 3529 5749 3581
rect 4485 3164 4491 3216
rect 4543 3164 4549 3216
rect 4910 3166 4916 3218
rect 4968 3166 4974 3218
rect 5307 3186 5335 3529
rect 5703 3186 5731 3529
rect 4493 2798 4541 3164
rect 4917 2798 4967 3166
rect 5289 3134 5295 3186
rect 5347 3134 5353 3186
rect 5685 3134 5691 3186
rect 5743 3134 5749 3186
rect 4485 2746 4491 2798
rect 4543 2746 4549 2798
rect 4910 2746 4916 2798
rect 4968 2746 4974 2798
rect 5307 2791 5335 3134
rect 5703 2791 5731 3134
rect 4493 2426 4541 2746
rect 4917 2428 4967 2746
rect 5289 2739 5295 2791
rect 5347 2739 5353 2791
rect 5685 2739 5691 2791
rect 5743 2739 5749 2791
rect 4485 2374 4491 2426
rect 4543 2374 4549 2426
rect 4910 2376 4916 2428
rect 4968 2376 4974 2428
rect 5307 2396 5335 2739
rect 5703 2396 5731 2739
rect 4493 2008 4541 2374
rect 4917 2008 4967 2376
rect 5289 2344 5295 2396
rect 5347 2344 5353 2396
rect 5685 2344 5691 2396
rect 5743 2344 5749 2396
rect 4485 1956 4491 2008
rect 4543 1956 4549 2008
rect 4910 1956 4916 2008
rect 4968 1956 4974 2008
rect 5307 2001 5335 2344
rect 5703 2001 5731 2344
rect 4493 1636 4541 1956
rect 4917 1638 4967 1956
rect 5289 1949 5295 2001
rect 5347 1949 5353 2001
rect 5685 1949 5691 2001
rect 5743 1949 5749 2001
rect 4485 1584 4491 1636
rect 4543 1584 4549 1636
rect 4910 1586 4916 1638
rect 4968 1586 4974 1638
rect 5307 1606 5335 1949
rect 5703 1606 5731 1949
rect 4493 1218 4541 1584
rect 4917 1218 4967 1586
rect 5289 1554 5295 1606
rect 5347 1554 5353 1606
rect 5685 1554 5691 1606
rect 5743 1554 5749 1606
rect 4485 1166 4491 1218
rect 4543 1166 4549 1218
rect 4910 1166 4916 1218
rect 4968 1166 4974 1218
rect 5307 1211 5335 1554
rect 5703 1211 5731 1554
rect 4493 846 4541 1166
rect 4917 848 4967 1166
rect 5289 1159 5295 1211
rect 5347 1159 5353 1211
rect 5685 1159 5691 1211
rect 5743 1159 5749 1211
rect 4485 794 4491 846
rect 4543 794 4549 846
rect 4910 796 4916 848
rect 4968 796 4974 848
rect 5307 816 5335 1159
rect 5703 816 5731 1159
rect 4493 428 4541 794
rect 4917 428 4967 796
rect 5289 764 5295 816
rect 5347 764 5353 816
rect 5685 764 5691 816
rect 5743 764 5749 816
rect 4485 376 4491 428
rect 4543 376 4549 428
rect 4910 376 4916 428
rect 4968 376 4974 428
rect 5307 421 5335 764
rect 5703 421 5731 764
rect 4493 -2 4541 376
rect 4917 -4 4967 376
rect 5289 369 5295 421
rect 5347 369 5353 421
rect 5685 369 5691 421
rect 5743 369 5749 421
rect 5307 28 5335 369
rect 5703 28 5731 369
rect 3595 -32 3647 -26
<< via1 >>
rect 3501 3847 3553 3856
rect 3501 3813 3510 3847
rect 3510 3813 3544 3847
rect 3544 3813 3553 3847
rect 3501 3804 3553 3813
rect 3501 3297 3553 3306
rect 3501 3263 3510 3297
rect 3510 3263 3544 3297
rect 3544 3263 3553 3297
rect 3501 3254 3553 3263
rect 3501 3057 3553 3066
rect 3501 3023 3510 3057
rect 3510 3023 3544 3057
rect 3544 3023 3553 3057
rect 3501 3014 3553 3023
rect 3501 2507 3553 2516
rect 3501 2473 3510 2507
rect 3510 2473 3544 2507
rect 3544 2473 3553 2507
rect 3501 2464 3553 2473
rect 3501 1477 3553 1486
rect 3501 1443 3510 1477
rect 3510 1443 3544 1477
rect 3544 1443 3553 1477
rect 3501 1434 3553 1443
rect 3501 927 3553 936
rect 3501 893 3510 927
rect 3510 893 3544 927
rect 3544 893 3553 927
rect 3501 884 3553 893
rect 3501 687 3553 696
rect 3501 653 3510 687
rect 3510 653 3544 687
rect 3544 653 3553 687
rect 3501 644 3553 653
rect 4491 5906 4543 5958
rect 4916 5906 4968 5958
rect 5295 5899 5347 5951
rect 5691 5899 5743 5951
rect 4491 5534 4543 5586
rect 4916 5536 4968 5588
rect 5295 5504 5347 5556
rect 5691 5504 5743 5556
rect 4491 5116 4543 5168
rect 4916 5116 4968 5168
rect 5295 5109 5347 5161
rect 5691 5109 5743 5161
rect 4491 4744 4543 4796
rect 4916 4746 4968 4798
rect 5295 4714 5347 4766
rect 5691 4714 5743 4766
rect 4491 4326 4543 4378
rect 4916 4326 4968 4378
rect 5295 4319 5347 4371
rect 5691 4319 5743 4371
rect 4491 3954 4543 4006
rect 4916 3956 4968 4008
rect 5295 3924 5347 3976
rect 5691 3924 5743 3976
rect 4155 3529 4207 3581
rect 4491 3536 4543 3588
rect 4916 3536 4968 3588
rect 4075 3134 4127 3186
rect 3995 2739 4047 2791
rect 3915 2344 3967 2396
rect 3835 1159 3887 1211
rect 3755 764 3807 816
rect 3675 369 3727 421
rect 3501 137 3553 146
rect 3501 103 3510 137
rect 3510 103 3544 137
rect 3544 103 3553 137
rect 3501 94 3553 103
rect 3595 -26 3647 26
rect 5295 3529 5347 3581
rect 5691 3529 5743 3581
rect 4491 3164 4543 3216
rect 4916 3166 4968 3218
rect 5295 3134 5347 3186
rect 5691 3134 5743 3186
rect 4491 2746 4543 2798
rect 4916 2746 4968 2798
rect 5295 2739 5347 2791
rect 5691 2739 5743 2791
rect 4491 2374 4543 2426
rect 4916 2376 4968 2428
rect 5295 2344 5347 2396
rect 5691 2344 5743 2396
rect 4491 1956 4543 2008
rect 4916 1956 4968 2008
rect 5295 1949 5347 2001
rect 5691 1949 5743 2001
rect 4491 1584 4543 1636
rect 4916 1586 4968 1638
rect 5295 1554 5347 1606
rect 5691 1554 5743 1606
rect 4491 1166 4543 1218
rect 4916 1166 4968 1218
rect 5295 1159 5347 1211
rect 5691 1159 5743 1211
rect 4491 794 4543 846
rect 4916 796 4968 848
rect 5295 764 5347 816
rect 5691 764 5743 816
rect 4491 376 4543 428
rect 4916 376 4968 428
rect 5295 369 5347 421
rect 5691 369 5743 421
<< metal2 >>
rect 4489 5960 4545 5969
rect 4489 5895 4545 5904
rect 4914 5960 4970 5969
rect 4914 5895 4970 5904
rect 5293 5953 5349 5962
rect 5293 5888 5349 5897
rect 5689 5953 5745 5962
rect 5689 5888 5745 5897
rect 4489 5588 4545 5597
rect 4489 5523 4545 5532
rect 4914 5590 4970 5599
rect 4914 5525 4970 5534
rect 5293 5558 5349 5567
rect 5293 5493 5349 5502
rect 5689 5558 5745 5567
rect 5689 5493 5745 5502
rect 4489 5170 4545 5179
rect 4489 5105 4545 5114
rect 4914 5170 4970 5179
rect 4914 5105 4970 5114
rect 5293 5163 5349 5172
rect 5293 5098 5349 5107
rect 5689 5163 5745 5172
rect 5689 5098 5745 5107
rect 4489 4798 4545 4807
rect 4489 4733 4545 4742
rect 4914 4800 4970 4809
rect 4914 4735 4970 4744
rect 5293 4768 5349 4777
rect 5293 4703 5349 4712
rect 5689 4768 5745 4777
rect 5689 4703 5745 4712
rect 4489 4380 4545 4389
rect 4489 4315 4545 4324
rect 4914 4380 4970 4389
rect 4914 4315 4970 4324
rect 5293 4373 5349 4382
rect 5293 4308 5349 4317
rect 5689 4373 5745 4382
rect 5689 4308 5745 4317
rect 4489 4008 4545 4017
rect 4489 3943 4545 3952
rect 4914 4010 4970 4019
rect 4914 3945 4970 3954
rect 5293 3978 5349 3987
rect 5293 3913 5349 3922
rect 5689 3978 5745 3987
rect 5689 3913 5745 3922
rect 3501 3856 3553 3862
rect 3501 3798 3553 3804
rect 3513 3569 3541 3798
rect 4489 3590 4545 3599
rect 4149 3569 4155 3581
rect 3513 3541 4155 3569
rect 4149 3529 4155 3541
rect 4207 3529 4213 3581
rect 4489 3525 4545 3534
rect 4914 3590 4970 3599
rect 4914 3525 4970 3534
rect 5293 3583 5349 3592
rect 5293 3518 5349 3527
rect 5689 3583 5745 3592
rect 5689 3518 5745 3527
rect 3501 3306 3553 3312
rect 3501 3248 3553 3254
rect 3513 3174 3541 3248
rect 4489 3218 4545 3227
rect 4069 3174 4075 3186
rect 3513 3146 4075 3174
rect 4069 3134 4075 3146
rect 4127 3134 4133 3186
rect 4489 3153 4545 3162
rect 4914 3220 4970 3229
rect 4914 3155 4970 3164
rect 5293 3188 5349 3197
rect 5293 3123 5349 3132
rect 5689 3188 5745 3197
rect 5689 3123 5745 3132
rect 3501 3066 3553 3072
rect 3501 3008 3553 3014
rect 3513 2779 3541 3008
rect 4489 2800 4545 2809
rect 3989 2779 3995 2791
rect 3513 2751 3995 2779
rect 3989 2739 3995 2751
rect 4047 2739 4053 2791
rect 4489 2735 4545 2744
rect 4914 2800 4970 2809
rect 4914 2735 4970 2744
rect 5293 2793 5349 2802
rect 5293 2728 5349 2737
rect 5689 2793 5745 2802
rect 5689 2728 5745 2737
rect 3501 2516 3553 2522
rect 3501 2458 3553 2464
rect 3513 2384 3541 2458
rect 4489 2428 4545 2437
rect 3909 2384 3915 2396
rect 3513 2356 3915 2384
rect 3909 2344 3915 2356
rect 3967 2344 3973 2396
rect 4489 2363 4545 2372
rect 4914 2430 4970 2439
rect 4914 2365 4970 2374
rect 5293 2398 5349 2407
rect 5293 2333 5349 2342
rect 5689 2398 5745 2407
rect 5689 2333 5745 2342
rect 4489 2010 4545 2019
rect 4489 1945 4545 1954
rect 4914 2010 4970 2019
rect 4914 1945 4970 1954
rect 5293 2003 5349 2012
rect 5293 1938 5349 1947
rect 5689 2003 5745 2012
rect 5689 1938 5745 1947
rect 4489 1638 4545 1647
rect 4489 1573 4545 1582
rect 4914 1640 4970 1649
rect 4914 1575 4970 1584
rect 5293 1608 5349 1617
rect 5293 1543 5349 1552
rect 5689 1608 5745 1617
rect 5689 1543 5745 1552
rect 3501 1486 3553 1492
rect 3501 1428 3553 1434
rect 3513 1199 3541 1428
rect 4489 1220 4545 1229
rect 3829 1199 3835 1211
rect 3513 1171 3835 1199
rect 3829 1159 3835 1171
rect 3887 1159 3893 1211
rect 4489 1155 4545 1164
rect 4914 1220 4970 1229
rect 4914 1155 4970 1164
rect 5293 1213 5349 1222
rect 5293 1148 5349 1157
rect 5689 1213 5745 1222
rect 5689 1148 5745 1157
rect 3501 936 3553 942
rect 3501 878 3553 884
rect 3513 804 3541 878
rect 4489 848 4545 857
rect 3749 804 3755 816
rect 3513 776 3755 804
rect 3749 764 3755 776
rect 3807 764 3813 816
rect 4489 783 4545 792
rect 4914 850 4970 859
rect 4914 785 4970 794
rect 5293 818 5349 827
rect 5293 753 5349 762
rect 5689 818 5745 827
rect 5689 753 5745 762
rect 3501 696 3553 702
rect 3501 638 3553 644
rect 3513 409 3541 638
rect 4489 430 4545 439
rect 3669 409 3675 421
rect 3513 381 3675 409
rect 3669 369 3675 381
rect 3727 369 3733 421
rect 4489 365 4545 374
rect 4914 430 4970 439
rect 4914 365 4970 374
rect 5293 423 5349 432
rect 5293 358 5349 367
rect 5689 423 5745 432
rect 5689 358 5745 367
rect 3501 146 3553 152
rect 3501 88 3553 94
rect 3513 14 3541 88
rect 3589 14 3595 26
rect 3513 -14 3595 14
rect 3589 -26 3595 -14
rect 3647 -26 3653 26
<< via2 >>
rect 4489 5958 4545 5960
rect 4489 5906 4491 5958
rect 4491 5906 4543 5958
rect 4543 5906 4545 5958
rect 4489 5904 4545 5906
rect 4914 5958 4970 5960
rect 4914 5906 4916 5958
rect 4916 5906 4968 5958
rect 4968 5906 4970 5958
rect 4914 5904 4970 5906
rect 5293 5951 5349 5953
rect 5293 5899 5295 5951
rect 5295 5899 5347 5951
rect 5347 5899 5349 5951
rect 5293 5897 5349 5899
rect 5689 5951 5745 5953
rect 5689 5899 5691 5951
rect 5691 5899 5743 5951
rect 5743 5899 5745 5951
rect 5689 5897 5745 5899
rect 4489 5586 4545 5588
rect 4489 5534 4491 5586
rect 4491 5534 4543 5586
rect 4543 5534 4545 5586
rect 4489 5532 4545 5534
rect 4914 5588 4970 5590
rect 4914 5536 4916 5588
rect 4916 5536 4968 5588
rect 4968 5536 4970 5588
rect 4914 5534 4970 5536
rect 5293 5556 5349 5558
rect 5293 5504 5295 5556
rect 5295 5504 5347 5556
rect 5347 5504 5349 5556
rect 5293 5502 5349 5504
rect 5689 5556 5745 5558
rect 5689 5504 5691 5556
rect 5691 5504 5743 5556
rect 5743 5504 5745 5556
rect 5689 5502 5745 5504
rect 4489 5168 4545 5170
rect 4489 5116 4491 5168
rect 4491 5116 4543 5168
rect 4543 5116 4545 5168
rect 4489 5114 4545 5116
rect 4914 5168 4970 5170
rect 4914 5116 4916 5168
rect 4916 5116 4968 5168
rect 4968 5116 4970 5168
rect 4914 5114 4970 5116
rect 5293 5161 5349 5163
rect 5293 5109 5295 5161
rect 5295 5109 5347 5161
rect 5347 5109 5349 5161
rect 5293 5107 5349 5109
rect 5689 5161 5745 5163
rect 5689 5109 5691 5161
rect 5691 5109 5743 5161
rect 5743 5109 5745 5161
rect 5689 5107 5745 5109
rect 4489 4796 4545 4798
rect 4489 4744 4491 4796
rect 4491 4744 4543 4796
rect 4543 4744 4545 4796
rect 4489 4742 4545 4744
rect 4914 4798 4970 4800
rect 4914 4746 4916 4798
rect 4916 4746 4968 4798
rect 4968 4746 4970 4798
rect 4914 4744 4970 4746
rect 5293 4766 5349 4768
rect 5293 4714 5295 4766
rect 5295 4714 5347 4766
rect 5347 4714 5349 4766
rect 5293 4712 5349 4714
rect 5689 4766 5745 4768
rect 5689 4714 5691 4766
rect 5691 4714 5743 4766
rect 5743 4714 5745 4766
rect 5689 4712 5745 4714
rect 4489 4378 4545 4380
rect 4489 4326 4491 4378
rect 4491 4326 4543 4378
rect 4543 4326 4545 4378
rect 4489 4324 4545 4326
rect 4914 4378 4970 4380
rect 4914 4326 4916 4378
rect 4916 4326 4968 4378
rect 4968 4326 4970 4378
rect 4914 4324 4970 4326
rect 5293 4371 5349 4373
rect 5293 4319 5295 4371
rect 5295 4319 5347 4371
rect 5347 4319 5349 4371
rect 5293 4317 5349 4319
rect 5689 4371 5745 4373
rect 5689 4319 5691 4371
rect 5691 4319 5743 4371
rect 5743 4319 5745 4371
rect 5689 4317 5745 4319
rect 4489 4006 4545 4008
rect 4489 3954 4491 4006
rect 4491 3954 4543 4006
rect 4543 3954 4545 4006
rect 4489 3952 4545 3954
rect 4914 4008 4970 4010
rect 4914 3956 4916 4008
rect 4916 3956 4968 4008
rect 4968 3956 4970 4008
rect 4914 3954 4970 3956
rect 5293 3976 5349 3978
rect 5293 3924 5295 3976
rect 5295 3924 5347 3976
rect 5347 3924 5349 3976
rect 5293 3922 5349 3924
rect 5689 3976 5745 3978
rect 5689 3924 5691 3976
rect 5691 3924 5743 3976
rect 5743 3924 5745 3976
rect 5689 3922 5745 3924
rect 4489 3588 4545 3590
rect 4489 3536 4491 3588
rect 4491 3536 4543 3588
rect 4543 3536 4545 3588
rect 4489 3534 4545 3536
rect 4914 3588 4970 3590
rect 4914 3536 4916 3588
rect 4916 3536 4968 3588
rect 4968 3536 4970 3588
rect 4914 3534 4970 3536
rect 5293 3581 5349 3583
rect 5293 3529 5295 3581
rect 5295 3529 5347 3581
rect 5347 3529 5349 3581
rect 5293 3527 5349 3529
rect 5689 3581 5745 3583
rect 5689 3529 5691 3581
rect 5691 3529 5743 3581
rect 5743 3529 5745 3581
rect 5689 3527 5745 3529
rect 4489 3216 4545 3218
rect 4489 3164 4491 3216
rect 4491 3164 4543 3216
rect 4543 3164 4545 3216
rect 4489 3162 4545 3164
rect 4914 3218 4970 3220
rect 4914 3166 4916 3218
rect 4916 3166 4968 3218
rect 4968 3166 4970 3218
rect 4914 3164 4970 3166
rect 5293 3186 5349 3188
rect 5293 3134 5295 3186
rect 5295 3134 5347 3186
rect 5347 3134 5349 3186
rect 5293 3132 5349 3134
rect 5689 3186 5745 3188
rect 5689 3134 5691 3186
rect 5691 3134 5743 3186
rect 5743 3134 5745 3186
rect 5689 3132 5745 3134
rect 4489 2798 4545 2800
rect 4489 2746 4491 2798
rect 4491 2746 4543 2798
rect 4543 2746 4545 2798
rect 4489 2744 4545 2746
rect 4914 2798 4970 2800
rect 4914 2746 4916 2798
rect 4916 2746 4968 2798
rect 4968 2746 4970 2798
rect 4914 2744 4970 2746
rect 5293 2791 5349 2793
rect 5293 2739 5295 2791
rect 5295 2739 5347 2791
rect 5347 2739 5349 2791
rect 5293 2737 5349 2739
rect 5689 2791 5745 2793
rect 5689 2739 5691 2791
rect 5691 2739 5743 2791
rect 5743 2739 5745 2791
rect 5689 2737 5745 2739
rect 4489 2426 4545 2428
rect 4489 2374 4491 2426
rect 4491 2374 4543 2426
rect 4543 2374 4545 2426
rect 4489 2372 4545 2374
rect 4914 2428 4970 2430
rect 4914 2376 4916 2428
rect 4916 2376 4968 2428
rect 4968 2376 4970 2428
rect 4914 2374 4970 2376
rect 5293 2396 5349 2398
rect 5293 2344 5295 2396
rect 5295 2344 5347 2396
rect 5347 2344 5349 2396
rect 5293 2342 5349 2344
rect 5689 2396 5745 2398
rect 5689 2344 5691 2396
rect 5691 2344 5743 2396
rect 5743 2344 5745 2396
rect 5689 2342 5745 2344
rect 4489 2008 4545 2010
rect 4489 1956 4491 2008
rect 4491 1956 4543 2008
rect 4543 1956 4545 2008
rect 4489 1954 4545 1956
rect 4914 2008 4970 2010
rect 4914 1956 4916 2008
rect 4916 1956 4968 2008
rect 4968 1956 4970 2008
rect 4914 1954 4970 1956
rect 5293 2001 5349 2003
rect 5293 1949 5295 2001
rect 5295 1949 5347 2001
rect 5347 1949 5349 2001
rect 5293 1947 5349 1949
rect 5689 2001 5745 2003
rect 5689 1949 5691 2001
rect 5691 1949 5743 2001
rect 5743 1949 5745 2001
rect 5689 1947 5745 1949
rect 4489 1636 4545 1638
rect 4489 1584 4491 1636
rect 4491 1584 4543 1636
rect 4543 1584 4545 1636
rect 4489 1582 4545 1584
rect 4914 1638 4970 1640
rect 4914 1586 4916 1638
rect 4916 1586 4968 1638
rect 4968 1586 4970 1638
rect 4914 1584 4970 1586
rect 5293 1606 5349 1608
rect 5293 1554 5295 1606
rect 5295 1554 5347 1606
rect 5347 1554 5349 1606
rect 5293 1552 5349 1554
rect 5689 1606 5745 1608
rect 5689 1554 5691 1606
rect 5691 1554 5743 1606
rect 5743 1554 5745 1606
rect 5689 1552 5745 1554
rect 4489 1218 4545 1220
rect 4489 1166 4491 1218
rect 4491 1166 4543 1218
rect 4543 1166 4545 1218
rect 4489 1164 4545 1166
rect 4914 1218 4970 1220
rect 4914 1166 4916 1218
rect 4916 1166 4968 1218
rect 4968 1166 4970 1218
rect 4914 1164 4970 1166
rect 5293 1211 5349 1213
rect 5293 1159 5295 1211
rect 5295 1159 5347 1211
rect 5347 1159 5349 1211
rect 5293 1157 5349 1159
rect 5689 1211 5745 1213
rect 5689 1159 5691 1211
rect 5691 1159 5743 1211
rect 5743 1159 5745 1211
rect 5689 1157 5745 1159
rect 4489 846 4545 848
rect 4489 794 4491 846
rect 4491 794 4543 846
rect 4543 794 4545 846
rect 4489 792 4545 794
rect 4914 848 4970 850
rect 4914 796 4916 848
rect 4916 796 4968 848
rect 4968 796 4970 848
rect 4914 794 4970 796
rect 5293 816 5349 818
rect 5293 764 5295 816
rect 5295 764 5347 816
rect 5347 764 5349 816
rect 5293 762 5349 764
rect 5689 816 5745 818
rect 5689 764 5691 816
rect 5691 764 5743 816
rect 5743 764 5745 816
rect 5689 762 5745 764
rect 4489 428 4545 430
rect 4489 376 4491 428
rect 4491 376 4543 428
rect 4543 376 4545 428
rect 4489 374 4545 376
rect 4914 428 4970 430
rect 4914 376 4916 428
rect 4916 376 4968 428
rect 4968 376 4970 428
rect 4914 374 4970 376
rect 5293 421 5349 423
rect 5293 369 5295 421
rect 5295 369 5347 421
rect 5347 369 5349 421
rect 5293 367 5349 369
rect 5689 421 5745 423
rect 5689 369 5691 421
rect 5691 369 5743 421
rect 5743 369 5745 421
rect 5689 367 5745 369
<< metal3 >>
rect 4468 5960 4566 5981
rect 4468 5904 4489 5960
rect 4545 5904 4566 5960
rect 4468 5883 4566 5904
rect 4893 5960 4991 5981
rect 4893 5904 4914 5960
rect 4970 5904 4991 5960
rect 4893 5883 4991 5904
rect 5272 5953 5370 5974
rect 5272 5897 5293 5953
rect 5349 5897 5370 5953
rect 5272 5876 5370 5897
rect 5668 5953 5766 5974
rect 5668 5897 5689 5953
rect 5745 5897 5766 5953
rect 5668 5876 5766 5897
rect 4468 5588 4566 5609
rect 4468 5532 4489 5588
rect 4545 5532 4566 5588
rect 4468 5511 4566 5532
rect 4893 5590 4991 5611
rect 4893 5534 4914 5590
rect 4970 5534 4991 5590
rect 4893 5513 4991 5534
rect 5272 5558 5370 5579
rect 5272 5502 5293 5558
rect 5349 5502 5370 5558
rect 5272 5481 5370 5502
rect 5668 5558 5766 5579
rect 5668 5502 5689 5558
rect 5745 5502 5766 5558
rect 5668 5481 5766 5502
rect 4468 5170 4566 5191
rect 4468 5114 4489 5170
rect 4545 5114 4566 5170
rect 4468 5093 4566 5114
rect 4893 5170 4991 5191
rect 4893 5114 4914 5170
rect 4970 5114 4991 5170
rect 4893 5093 4991 5114
rect 5272 5163 5370 5184
rect 5272 5107 5293 5163
rect 5349 5107 5370 5163
rect 5272 5086 5370 5107
rect 5668 5163 5766 5184
rect 5668 5107 5689 5163
rect 5745 5107 5766 5163
rect 5668 5086 5766 5107
rect 4468 4798 4566 4819
rect 4468 4742 4489 4798
rect 4545 4742 4566 4798
rect 4468 4721 4566 4742
rect 4893 4800 4991 4821
rect 4893 4744 4914 4800
rect 4970 4744 4991 4800
rect 4893 4723 4991 4744
rect 5272 4768 5370 4789
rect 5272 4712 5293 4768
rect 5349 4712 5370 4768
rect 5272 4691 5370 4712
rect 5668 4768 5766 4789
rect 5668 4712 5689 4768
rect 5745 4712 5766 4768
rect 5668 4691 5766 4712
rect 4468 4380 4566 4401
rect 4468 4324 4489 4380
rect 4545 4324 4566 4380
rect 4468 4303 4566 4324
rect 4893 4380 4991 4401
rect 4893 4324 4914 4380
rect 4970 4324 4991 4380
rect 4893 4303 4991 4324
rect 5272 4373 5370 4394
rect 5272 4317 5293 4373
rect 5349 4317 5370 4373
rect 5272 4296 5370 4317
rect 5668 4373 5766 4394
rect 5668 4317 5689 4373
rect 5745 4317 5766 4373
rect 5668 4296 5766 4317
rect 4468 4008 4566 4029
rect 4468 3952 4489 4008
rect 4545 3952 4566 4008
rect 4468 3931 4566 3952
rect 4893 4010 4991 4031
rect 4893 3954 4914 4010
rect 4970 3954 4991 4010
rect 4893 3933 4991 3954
rect 5272 3978 5370 3999
rect 5272 3922 5293 3978
rect 5349 3922 5370 3978
rect 5272 3901 5370 3922
rect 5668 3978 5766 3999
rect 5668 3922 5689 3978
rect 5745 3922 5766 3978
rect 5668 3901 5766 3922
rect 2130 3513 2228 3611
rect 2555 3513 2653 3611
rect 2934 3506 3032 3604
rect 3330 3506 3428 3604
rect 4468 3590 4566 3611
rect 4468 3534 4489 3590
rect 4545 3534 4566 3590
rect 4468 3513 4566 3534
rect 4893 3590 4991 3611
rect 4893 3534 4914 3590
rect 4970 3534 4991 3590
rect 4893 3513 4991 3534
rect 5272 3583 5370 3604
rect 5272 3527 5293 3583
rect 5349 3527 5370 3583
rect 5272 3506 5370 3527
rect 5668 3583 5766 3604
rect 5668 3527 5689 3583
rect 5745 3527 5766 3583
rect 5668 3506 5766 3527
rect 4468 3218 4566 3239
rect 4468 3162 4489 3218
rect 4545 3162 4566 3218
rect 4468 3141 4566 3162
rect 4893 3220 4991 3241
rect 4893 3164 4914 3220
rect 4970 3164 4991 3220
rect 4893 3143 4991 3164
rect 5272 3188 5370 3209
rect 5272 3132 5293 3188
rect 5349 3132 5370 3188
rect 5272 3111 5370 3132
rect 5668 3188 5766 3209
rect 5668 3132 5689 3188
rect 5745 3132 5766 3188
rect 5668 3111 5766 3132
rect 836 2716 934 2814
rect 1232 2716 1330 2814
rect 2130 2723 2228 2821
rect 2555 2723 2653 2821
rect 2934 2716 3032 2814
rect 3330 2716 3428 2814
rect 4468 2800 4566 2821
rect 4468 2744 4489 2800
rect 4545 2744 4566 2800
rect 4468 2723 4566 2744
rect 4893 2800 4991 2821
rect 4893 2744 4914 2800
rect 4970 2744 4991 2800
rect 4893 2723 4991 2744
rect 5272 2793 5370 2814
rect 5272 2737 5293 2793
rect 5349 2737 5370 2793
rect 5272 2716 5370 2737
rect 5668 2793 5766 2814
rect 5668 2737 5689 2793
rect 5745 2737 5766 2793
rect 5668 2716 5766 2737
rect 4468 2428 4566 2449
rect 4468 2372 4489 2428
rect 4545 2372 4566 2428
rect 4468 2351 4566 2372
rect 4893 2430 4991 2451
rect 4893 2374 4914 2430
rect 4970 2374 4991 2430
rect 4893 2353 4991 2374
rect 5272 2398 5370 2419
rect 5272 2342 5293 2398
rect 5349 2342 5370 2398
rect 5272 2321 5370 2342
rect 5668 2398 5766 2419
rect 5668 2342 5689 2398
rect 5745 2342 5766 2398
rect 5668 2321 5766 2342
rect 4468 2010 4566 2031
rect 4468 1954 4489 2010
rect 4545 1954 4566 2010
rect 4468 1933 4566 1954
rect 4893 2010 4991 2031
rect 4893 1954 4914 2010
rect 4970 1954 4991 2010
rect 4893 1933 4991 1954
rect 5272 2003 5370 2024
rect 5272 1947 5293 2003
rect 5349 1947 5370 2003
rect 5272 1926 5370 1947
rect 5668 2003 5766 2024
rect 5668 1947 5689 2003
rect 5745 1947 5766 2003
rect 5668 1926 5766 1947
rect 4468 1638 4566 1659
rect 4468 1582 4489 1638
rect 4545 1582 4566 1638
rect 4468 1561 4566 1582
rect 4893 1640 4991 1661
rect 4893 1584 4914 1640
rect 4970 1584 4991 1640
rect 4893 1563 4991 1584
rect 5272 1608 5370 1629
rect 5272 1552 5293 1608
rect 5349 1552 5370 1608
rect 5272 1531 5370 1552
rect 5668 1608 5766 1629
rect 5668 1552 5689 1608
rect 5745 1552 5766 1608
rect 5668 1531 5766 1552
rect 2130 1143 2228 1241
rect 2555 1143 2653 1241
rect 2934 1136 3032 1234
rect 3330 1136 3428 1234
rect 4468 1220 4566 1241
rect 4468 1164 4489 1220
rect 4545 1164 4566 1220
rect 4468 1143 4566 1164
rect 4893 1220 4991 1241
rect 4893 1164 4914 1220
rect 4970 1164 4991 1220
rect 4893 1143 4991 1164
rect 5272 1213 5370 1234
rect 5272 1157 5293 1213
rect 5349 1157 5370 1213
rect 5272 1136 5370 1157
rect 5668 1213 5766 1234
rect 5668 1157 5689 1213
rect 5745 1157 5766 1213
rect 5668 1136 5766 1157
rect 4468 848 4566 869
rect 4468 792 4489 848
rect 4545 792 4566 848
rect 4468 771 4566 792
rect 4893 850 4991 871
rect 4893 794 4914 850
rect 4970 794 4991 850
rect 4893 773 4991 794
rect 5272 818 5370 839
rect 5272 762 5293 818
rect 5349 762 5370 818
rect 5272 741 5370 762
rect 5668 818 5766 839
rect 5668 762 5689 818
rect 5745 762 5766 818
rect 5668 741 5766 762
rect 836 346 934 444
rect 1232 346 1330 444
rect 2130 353 2228 451
rect 2555 353 2653 451
rect 2934 346 3032 444
rect 3330 346 3428 444
rect 4468 430 4566 451
rect 4468 374 4489 430
rect 4545 374 4566 430
rect 4468 353 4566 374
rect 4893 430 4991 451
rect 4893 374 4914 430
rect 4970 374 4991 430
rect 4893 353 4991 374
rect 5272 423 5370 444
rect 5272 367 5293 423
rect 5349 367 5370 423
rect 5272 346 5370 367
rect 5668 423 5766 444
rect 5668 367 5689 423
rect 5745 367 5766 423
rect 5668 346 5766 367
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 5288 0 1 5888
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 5289 0 1 5893
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 4484 0 1 5895
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 4485 0 1 5900
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 5288 0 1 5493
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 5289 0 1 5498
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 4484 0 1 5523
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 4485 0 1 5528
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 5288 0 1 5098
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 5289 0 1 5103
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 4484 0 1 5105
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 4485 0 1 5110
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 5288 0 1 4703
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 5289 0 1 4708
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 4484 0 1 4733
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 4485 0 1 4738
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 5288 0 1 4308
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 5289 0 1 4313
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 4484 0 1 4315
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 4485 0 1 4320
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 5288 0 1 3913
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 5289 0 1 3918
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 4484 0 1 3943
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 4485 0 1 3948
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 5288 0 1 3518
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 5289 0 1 3523
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 4484 0 1 3525
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 4485 0 1 3530
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 5288 0 1 3123
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 5289 0 1 3128
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 4484 0 1 3153
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 4485 0 1 3158
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 5288 0 1 2728
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1634918361
transform 1 0 5289 0 1 2733
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1634918361
transform 1 0 4484 0 1 2735
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1634918361
transform 1 0 4485 0 1 2740
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1634918361
transform 1 0 5288 0 1 2333
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1634918361
transform 1 0 5289 0 1 2338
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1634918361
transform 1 0 4484 0 1 2363
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1634918361
transform 1 0 4485 0 1 2368
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1634918361
transform 1 0 5288 0 1 1938
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1634918361
transform 1 0 5289 0 1 1943
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1634918361
transform 1 0 4484 0 1 1945
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1634918361
transform 1 0 4485 0 1 1950
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1634918361
transform 1 0 5288 0 1 1543
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1634918361
transform 1 0 5289 0 1 1548
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1634918361
transform 1 0 4484 0 1 1573
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1634918361
transform 1 0 4485 0 1 1578
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1634918361
transform 1 0 5288 0 1 1148
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1634918361
transform 1 0 5289 0 1 1153
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1634918361
transform 1 0 4484 0 1 1155
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1634918361
transform 1 0 4485 0 1 1160
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1634918361
transform 1 0 5288 0 1 753
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1634918361
transform 1 0 5289 0 1 758
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1634918361
transform 1 0 4484 0 1 783
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1634918361
transform 1 0 4485 0 1 788
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1634918361
transform 1 0 5288 0 1 358
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1634918361
transform 1 0 5289 0 1 363
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1634918361
transform 1 0 4484 0 1 365
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1634918361
transform 1 0 4485 0 1 370
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1634918361
transform 1 0 4909 0 1 5895
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1634918361
transform 1 0 4910 0 1 5900
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1634918361
transform 1 0 5684 0 1 5888
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1634918361
transform 1 0 5685 0 1 5893
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1634918361
transform 1 0 4909 0 1 5525
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1634918361
transform 1 0 4910 0 1 5530
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1634918361
transform 1 0 5684 0 1 5493
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1634918361
transform 1 0 5685 0 1 5498
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1634918361
transform 1 0 4909 0 1 5105
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1634918361
transform 1 0 4910 0 1 5110
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1634918361
transform 1 0 5684 0 1 5098
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1634918361
transform 1 0 5685 0 1 5103
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1634918361
transform 1 0 4909 0 1 4735
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1634918361
transform 1 0 4910 0 1 4740
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1634918361
transform 1 0 5684 0 1 4703
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1634918361
transform 1 0 5685 0 1 4708
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1634918361
transform 1 0 4909 0 1 4315
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1634918361
transform 1 0 4910 0 1 4320
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1634918361
transform 1 0 5684 0 1 4308
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1634918361
transform 1 0 5685 0 1 4313
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1634918361
transform 1 0 4909 0 1 3945
box 0 0 1 1
use contact_19  contact_19_40
timestamp 1634918361
transform 1 0 4910 0 1 3950
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1634918361
transform 1 0 5684 0 1 3913
box 0 0 1 1
use contact_19  contact_19_41
timestamp 1634918361
transform 1 0 5685 0 1 3918
box 0 0 1 1
use contact_7  contact_7_42
timestamp 1634918361
transform 1 0 4909 0 1 3525
box 0 0 1 1
use contact_19  contact_19_42
timestamp 1634918361
transform 1 0 4910 0 1 3530
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1634918361
transform 1 0 5684 0 1 3518
box 0 0 1 1
use contact_19  contact_19_43
timestamp 1634918361
transform 1 0 5685 0 1 3523
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1634918361
transform 1 0 4909 0 1 3155
box 0 0 1 1
use contact_19  contact_19_44
timestamp 1634918361
transform 1 0 4910 0 1 3160
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1634918361
transform 1 0 5684 0 1 3123
box 0 0 1 1
use contact_19  contact_19_45
timestamp 1634918361
transform 1 0 5685 0 1 3128
box 0 0 1 1
use contact_7  contact_7_46
timestamp 1634918361
transform 1 0 4909 0 1 2735
box 0 0 1 1
use contact_19  contact_19_46
timestamp 1634918361
transform 1 0 4910 0 1 2740
box 0 0 1 1
use contact_7  contact_7_47
timestamp 1634918361
transform 1 0 5684 0 1 2728
box 0 0 1 1
use contact_19  contact_19_47
timestamp 1634918361
transform 1 0 5685 0 1 2733
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1634918361
transform 1 0 4909 0 1 2365
box 0 0 1 1
use contact_19  contact_19_48
timestamp 1634918361
transform 1 0 4910 0 1 2370
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1634918361
transform 1 0 5684 0 1 2333
box 0 0 1 1
use contact_19  contact_19_49
timestamp 1634918361
transform 1 0 5685 0 1 2338
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1634918361
transform 1 0 4909 0 1 1945
box 0 0 1 1
use contact_19  contact_19_50
timestamp 1634918361
transform 1 0 4910 0 1 1950
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1634918361
transform 1 0 5684 0 1 1938
box 0 0 1 1
use contact_19  contact_19_51
timestamp 1634918361
transform 1 0 5685 0 1 1943
box 0 0 1 1
use contact_7  contact_7_52
timestamp 1634918361
transform 1 0 4909 0 1 1575
box 0 0 1 1
use contact_19  contact_19_52
timestamp 1634918361
transform 1 0 4910 0 1 1580
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1634918361
transform 1 0 5684 0 1 1543
box 0 0 1 1
use contact_19  contact_19_53
timestamp 1634918361
transform 1 0 5685 0 1 1548
box 0 0 1 1
use contact_7  contact_7_54
timestamp 1634918361
transform 1 0 4909 0 1 1155
box 0 0 1 1
use contact_19  contact_19_54
timestamp 1634918361
transform 1 0 4910 0 1 1160
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1634918361
transform 1 0 5684 0 1 1148
box 0 0 1 1
use contact_19  contact_19_55
timestamp 1634918361
transform 1 0 5685 0 1 1153
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1634918361
transform 1 0 4909 0 1 785
box 0 0 1 1
use contact_19  contact_19_56
timestamp 1634918361
transform 1 0 4910 0 1 790
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1634918361
transform 1 0 5684 0 1 753
box 0 0 1 1
use contact_19  contact_19_57
timestamp 1634918361
transform 1 0 5685 0 1 758
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1634918361
transform 1 0 4909 0 1 365
box 0 0 1 1
use contact_19  contact_19_58
timestamp 1634918361
transform 1 0 4910 0 1 370
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1634918361
transform 1 0 5684 0 1 358
box 0 0 1 1
use contact_19  contact_19_59
timestamp 1634918361
transform 1 0 5685 0 1 363
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1634918361
transform 1 0 4149 0 1 3523
box 0 0 1 1
use contact_19  contact_19_60
timestamp 1634918361
transform 1 0 3495 0 1 3798
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 3498 0 1 3797
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1634918361
transform 1 0 4069 0 1 3128
box 0 0 1 1
use contact_19  contact_19_61
timestamp 1634918361
transform 1 0 3495 0 1 3248
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 3498 0 1 3247
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1634918361
transform 1 0 3989 0 1 2733
box 0 0 1 1
use contact_19  contact_19_62
timestamp 1634918361
transform 1 0 3495 0 1 3008
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 3498 0 1 3007
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1634918361
transform 1 0 3909 0 1 2338
box 0 0 1 1
use contact_19  contact_19_63
timestamp 1634918361
transform 1 0 3495 0 1 2458
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 3498 0 1 2457
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1634918361
transform 1 0 3829 0 1 1153
box 0 0 1 1
use contact_19  contact_19_64
timestamp 1634918361
transform 1 0 3495 0 1 1428
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 3498 0 1 1427
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1634918361
transform 1 0 3749 0 1 758
box 0 0 1 1
use contact_19  contact_19_65
timestamp 1634918361
transform 1 0 3495 0 1 878
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 3498 0 1 877
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1634918361
transform 1 0 3669 0 1 363
box 0 0 1 1
use contact_19  contact_19_66
timestamp 1634918361
transform 1 0 3495 0 1 638
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 3498 0 1 637
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1634918361
transform 1 0 3589 0 1 -32
box 0 0 1 1
use contact_19  contact_19_67
timestamp 1634918361
transform 1 0 3495 0 1 88
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 3498 0 1 87
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1634918361
transform 1 0 4148 0 1 6100
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1634918361
transform 1 0 3828 0 1 5992
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1634918361
transform 1 0 4148 0 1 5692
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1634918361
transform 1 0 3748 0 1 5800
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1634918361
transform 1 0 4148 0 1 5310
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1634918361
transform 1 0 3668 0 1 5202
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1634918361
transform 1 0 4148 0 1 4902
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1634918361
transform 1 0 3588 0 1 5010
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1634918361
transform 1 0 4068 0 1 4520
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1634918361
transform 1 0 3828 0 1 4412
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1634918361
transform 1 0 4068 0 1 4112
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1634918361
transform 1 0 3748 0 1 4220
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1634918361
transform 1 0 4068 0 1 3730
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1634918361
transform 1 0 3668 0 1 3622
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1634918361
transform 1 0 4068 0 1 3322
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1634918361
transform 1 0 3588 0 1 3430
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1634918361
transform 1 0 3988 0 1 2940
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1634918361
transform 1 0 3828 0 1 2832
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1634918361
transform 1 0 3988 0 1 2532
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1634918361
transform 1 0 3748 0 1 2640
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1634918361
transform 1 0 3988 0 1 2150
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1634918361
transform 1 0 3668 0 1 2042
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1634918361
transform 1 0 3988 0 1 1742
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1634918361
transform 1 0 3588 0 1 1850
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1634918361
transform 1 0 3908 0 1 1360
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1634918361
transform 1 0 3828 0 1 1252
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1634918361
transform 1 0 3908 0 1 952
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1634918361
transform 1 0 3748 0 1 1060
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1634918361
transform 1 0 3908 0 1 570
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1634918361
transform 1 0 3668 0 1 462
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1634918361
transform 1 0 3908 0 1 162
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1634918361
transform 1 0 3588 0 1 270
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1634918361
transform 1 0 240 0 1 2961
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 512 0 1 2957
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1634918361
transform 1 0 160 0 1 2511
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 432 0 1 2507
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1634918361
transform 1 0 80 0 1 591
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 512 0 1 587
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1634918361
transform 1 0 0 0 1 141
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 432 0 1 137
box 0 0 1 1
use and2_dec  and2_dec_0
timestamp 1634918361
transform 1 0 4247 0 -1 6320
box 70 -56 1636 490
use and2_dec  and2_dec_1
timestamp 1634918361
transform 1 0 4247 0 1 5530
box 70 -56 1636 490
use and2_dec  and2_dec_2
timestamp 1634918361
transform 1 0 4247 0 -1 5530
box 70 -56 1636 490
use and2_dec  and2_dec_3
timestamp 1634918361
transform 1 0 4247 0 1 4740
box 70 -56 1636 490
use and2_dec  and2_dec_4
timestamp 1634918361
transform 1 0 4247 0 -1 4740
box 70 -56 1636 490
use and2_dec  and2_dec_5
timestamp 1634918361
transform 1 0 4247 0 1 3950
box 70 -56 1636 490
use and2_dec  and2_dec_6
timestamp 1634918361
transform 1 0 4247 0 -1 3950
box 70 -56 1636 490
use and2_dec  and2_dec_7
timestamp 1634918361
transform 1 0 4247 0 1 3160
box 70 -56 1636 490
use and2_dec  and2_dec_8
timestamp 1634918361
transform 1 0 4247 0 -1 3160
box 70 -56 1636 490
use and2_dec  and2_dec_9
timestamp 1634918361
transform 1 0 4247 0 1 2370
box 70 -56 1636 490
use and2_dec  and2_dec_10
timestamp 1634918361
transform 1 0 4247 0 -1 2370
box 70 -56 1636 490
use and2_dec  and2_dec_11
timestamp 1634918361
transform 1 0 4247 0 1 1580
box 70 -56 1636 490
use and2_dec  and2_dec_12
timestamp 1634918361
transform 1 0 4247 0 -1 1580
box 70 -56 1636 490
use and2_dec  and2_dec_13
timestamp 1634918361
transform 1 0 4247 0 1 790
box 70 -56 1636 490
use and2_dec  and2_dec_14
timestamp 1634918361
transform 1 0 4247 0 -1 790
box 70 -56 1636 490
use and2_dec  and2_dec_15
timestamp 1634918361
transform 1 0 4247 0 1 0
box 70 -56 1636 490
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1634918361
transform 1 0 367 0 1 2370
box 61 -56 3178 1636
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1634918361
transform 1 0 367 0 1 0
box 61 -56 3178 1636
<< labels >>
rlabel metal1 s 19 0 47 3950 4 addr_0
port 1 nsew
rlabel metal1 s 99 0 127 3950 4 addr_1
port 2 nsew
rlabel metal1 s 179 0 207 3950 4 addr_2
port 3 nsew
rlabel metal1 s 259 0 287 3950 4 addr_3
port 4 nsew
rlabel locali s 5576 120 5576 120 4 decode_0
port 5 nsew
rlabel locali s 5576 670 5576 670 4 decode_1
port 6 nsew
rlabel locali s 5576 910 5576 910 4 decode_2
port 7 nsew
rlabel locali s 5576 1460 5576 1460 4 decode_3
port 8 nsew
rlabel locali s 5576 1700 5576 1700 4 decode_4
port 9 nsew
rlabel locali s 5576 2250 5576 2250 4 decode_5
port 10 nsew
rlabel locali s 5576 2490 5576 2490 4 decode_6
port 11 nsew
rlabel locali s 5576 3040 5576 3040 4 decode_7
port 12 nsew
rlabel locali s 5576 3280 5576 3280 4 decode_8
port 13 nsew
rlabel locali s 5576 3830 5576 3830 4 decode_9
port 14 nsew
rlabel locali s 5576 4070 5576 4070 4 decode_10
port 15 nsew
rlabel locali s 5576 4620 5576 4620 4 decode_11
port 16 nsew
rlabel locali s 5576 4860 5576 4860 4 decode_12
port 17 nsew
rlabel locali s 5576 5410 5576 5410 4 decode_13
port 18 nsew
rlabel locali s 5576 5650 5576 5650 4 decode_14
port 19 nsew
rlabel locali s 5576 6200 5576 6200 4 decode_15
port 20 nsew
rlabel metal1 s 3607 0 3635 6348 4 predecode_0
port 21 nsew
rlabel metal1 s 3687 0 3715 6348 4 predecode_1
port 22 nsew
rlabel metal1 s 3767 0 3795 6348 4 predecode_2
port 23 nsew
rlabel metal1 s 3847 0 3875 6348 4 predecode_3
port 24 nsew
rlabel metal1 s 3927 0 3955 6348 4 predecode_4
port 25 nsew
rlabel metal1 s 4007 0 4035 6348 4 predecode_5
port 26 nsew
rlabel metal1 s 4087 0 4115 6348 4 predecode_6
port 27 nsew
rlabel metal1 s 4167 0 4195 6348 4 predecode_7
port 28 nsew
rlabel metal3 s 5668 1926 5766 2024 4 vdd
port 29 nsew
rlabel metal3 s 4893 2723 4991 2821 4 vdd
port 29 nsew
rlabel metal3 s 3330 346 3428 444 4 vdd
port 29 nsew
rlabel metal3 s 5668 4296 5766 4394 4 vdd
port 29 nsew
rlabel metal3 s 5668 2321 5766 2419 4 vdd
port 29 nsew
rlabel metal3 s 4893 3513 4991 3611 4 vdd
port 29 nsew
rlabel metal3 s 4893 4303 4991 4401 4 vdd
port 29 nsew
rlabel metal3 s 4893 1933 4991 2031 4 vdd
port 29 nsew
rlabel metal3 s 4893 5513 4991 5611 4 vdd
port 29 nsew
rlabel metal3 s 4893 3933 4991 4031 4 vdd
port 29 nsew
rlabel metal3 s 1232 346 1330 444 4 vdd
port 29 nsew
rlabel metal3 s 5668 5481 5766 5579 4 vdd
port 29 nsew
rlabel metal3 s 5668 346 5766 444 4 vdd
port 29 nsew
rlabel metal3 s 5668 3111 5766 3209 4 vdd
port 29 nsew
rlabel metal3 s 2555 1143 2653 1241 4 vdd
port 29 nsew
rlabel metal3 s 5668 2716 5766 2814 4 vdd
port 29 nsew
rlabel metal3 s 5668 4691 5766 4789 4 vdd
port 29 nsew
rlabel metal3 s 2555 2723 2653 2821 4 vdd
port 29 nsew
rlabel metal3 s 3330 1136 3428 1234 4 vdd
port 29 nsew
rlabel metal3 s 4893 3143 4991 3241 4 vdd
port 29 nsew
rlabel metal3 s 4893 5883 4991 5981 4 vdd
port 29 nsew
rlabel metal3 s 2555 3513 2653 3611 4 vdd
port 29 nsew
rlabel metal3 s 1232 2716 1330 2814 4 vdd
port 29 nsew
rlabel metal3 s 4893 1563 4991 1661 4 vdd
port 29 nsew
rlabel metal3 s 5668 1136 5766 1234 4 vdd
port 29 nsew
rlabel metal3 s 4893 353 4991 451 4 vdd
port 29 nsew
rlabel metal3 s 5668 3901 5766 3999 4 vdd
port 29 nsew
rlabel metal3 s 5668 5086 5766 5184 4 vdd
port 29 nsew
rlabel metal3 s 4893 2353 4991 2451 4 vdd
port 29 nsew
rlabel metal3 s 5668 5876 5766 5974 4 vdd
port 29 nsew
rlabel metal3 s 4893 773 4991 871 4 vdd
port 29 nsew
rlabel metal3 s 5668 3506 5766 3604 4 vdd
port 29 nsew
rlabel metal3 s 3330 3506 3428 3604 4 vdd
port 29 nsew
rlabel metal3 s 5668 741 5766 839 4 vdd
port 29 nsew
rlabel metal3 s 5668 1531 5766 1629 4 vdd
port 29 nsew
rlabel metal3 s 4893 4723 4991 4821 4 vdd
port 29 nsew
rlabel metal3 s 2555 353 2653 451 4 vdd
port 29 nsew
rlabel metal3 s 3330 2716 3428 2814 4 vdd
port 29 nsew
rlabel metal3 s 4893 5093 4991 5191 4 vdd
port 29 nsew
rlabel metal3 s 4893 1143 4991 1241 4 vdd
port 29 nsew
rlabel metal3 s 4468 1933 4566 2031 4 gnd
port 30 nsew
rlabel metal3 s 2934 3506 3032 3604 4 gnd
port 30 nsew
rlabel metal3 s 2934 346 3032 444 4 gnd
port 30 nsew
rlabel metal3 s 4468 3931 4566 4029 4 gnd
port 30 nsew
rlabel metal3 s 5272 4691 5370 4789 4 gnd
port 30 nsew
rlabel metal3 s 4468 4303 4566 4401 4 gnd
port 30 nsew
rlabel metal3 s 5272 3901 5370 3999 4 gnd
port 30 nsew
rlabel metal3 s 4468 353 4566 451 4 gnd
port 30 nsew
rlabel metal3 s 4468 771 4566 869 4 gnd
port 30 nsew
rlabel metal3 s 4468 1143 4566 1241 4 gnd
port 30 nsew
rlabel metal3 s 5272 3111 5370 3209 4 gnd
port 30 nsew
rlabel metal3 s 5272 1926 5370 2024 4 gnd
port 30 nsew
rlabel metal3 s 4468 5883 4566 5981 4 gnd
port 30 nsew
rlabel metal3 s 2130 2723 2228 2821 4 gnd
port 30 nsew
rlabel metal3 s 5272 1136 5370 1234 4 gnd
port 30 nsew
rlabel metal3 s 4468 3513 4566 3611 4 gnd
port 30 nsew
rlabel metal3 s 4468 2723 4566 2821 4 gnd
port 30 nsew
rlabel metal3 s 836 2716 934 2814 4 gnd
port 30 nsew
rlabel metal3 s 5272 2716 5370 2814 4 gnd
port 30 nsew
rlabel metal3 s 4468 1561 4566 1659 4 gnd
port 30 nsew
rlabel metal3 s 2130 3513 2228 3611 4 gnd
port 30 nsew
rlabel metal3 s 5272 5086 5370 5184 4 gnd
port 30 nsew
rlabel metal3 s 4468 5093 4566 5191 4 gnd
port 30 nsew
rlabel metal3 s 5272 5481 5370 5579 4 gnd
port 30 nsew
rlabel metal3 s 4468 4721 4566 4819 4 gnd
port 30 nsew
rlabel metal3 s 4468 3141 4566 3239 4 gnd
port 30 nsew
rlabel metal3 s 2130 1143 2228 1241 4 gnd
port 30 nsew
rlabel metal3 s 5272 3506 5370 3604 4 gnd
port 30 nsew
rlabel metal3 s 5272 1531 5370 1629 4 gnd
port 30 nsew
rlabel metal3 s 2130 353 2228 451 4 gnd
port 30 nsew
rlabel metal3 s 836 346 934 444 4 gnd
port 30 nsew
rlabel metal3 s 2934 2716 3032 2814 4 gnd
port 30 nsew
rlabel metal3 s 5272 4296 5370 4394 4 gnd
port 30 nsew
rlabel metal3 s 5272 2321 5370 2419 4 gnd
port 30 nsew
rlabel metal3 s 4468 2351 4566 2449 4 gnd
port 30 nsew
rlabel metal3 s 4468 5511 4566 5609 4 gnd
port 30 nsew
rlabel metal3 s 5272 5876 5370 5974 4 gnd
port 30 nsew
rlabel metal3 s 5272 346 5370 444 4 gnd
port 30 nsew
rlabel metal3 s 2934 1136 3032 1234 4 gnd
port 30 nsew
rlabel metal3 s 5272 741 5370 839 4 gnd
port 30 nsew
<< properties >>
string FIXED_BBOX 3589 -32 3653 0
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 975206
string GDS_START 938582
<< end >>
