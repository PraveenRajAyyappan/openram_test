magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1260 -1260 25562 19956
<< locali >>
rect 16089 14445 16123 14461
rect 16123 14411 16269 14445
rect 16089 14395 16123 14411
rect 8095 14205 8129 14221
rect 7949 14171 8095 14205
rect 8095 14155 8129 14171
rect 16089 14205 16123 14221
rect 16123 14171 16269 14205
rect 16089 14155 16123 14171
rect 8095 13655 8129 13671
rect 7949 13621 8095 13655
rect 8095 13605 8129 13621
rect 16089 13655 16123 13671
rect 16123 13621 16269 13655
rect 16089 13605 16123 13621
rect 8095 13415 8129 13431
rect 7949 13381 8095 13415
rect 8095 13365 8129 13381
rect 16089 13415 16123 13431
rect 16123 13381 16269 13415
rect 16089 13365 16123 13381
rect 8095 12865 8129 12881
rect 7949 12831 8095 12865
rect 8095 12815 8129 12831
rect 16089 12865 16123 12881
rect 16123 12831 16269 12865
rect 16089 12815 16123 12831
rect 8095 12625 8129 12641
rect 7949 12591 8095 12625
rect 8095 12575 8129 12591
rect 16089 12625 16123 12641
rect 16123 12591 16269 12625
rect 16089 12575 16123 12591
rect 8095 12075 8129 12091
rect 7949 12041 8095 12075
rect 8095 12025 8129 12041
rect 16089 12075 16123 12091
rect 16123 12041 16269 12075
rect 16089 12025 16123 12041
rect 8095 11835 8129 11851
rect 7949 11801 8095 11835
rect 8095 11785 8129 11801
rect 16089 11835 16123 11851
rect 16123 11801 16269 11835
rect 16089 11785 16123 11801
rect 8095 11285 8129 11301
rect 7949 11251 8095 11285
rect 8095 11235 8129 11251
rect 16089 11285 16123 11301
rect 16123 11251 16269 11285
rect 16089 11235 16123 11251
rect 8095 11045 8129 11061
rect 7949 11011 8095 11045
rect 8095 10995 8129 11011
rect 16089 11045 16123 11061
rect 16123 11011 16269 11045
rect 16089 10995 16123 11011
rect 8095 10495 8129 10511
rect 7949 10461 8095 10495
rect 8095 10445 8129 10461
rect 16089 10495 16123 10511
rect 16123 10461 16269 10495
rect 16089 10445 16123 10461
rect 8095 10255 8129 10271
rect 7949 10221 8095 10255
rect 8095 10205 8129 10221
rect 16089 10255 16123 10271
rect 16123 10221 16269 10255
rect 16089 10205 16123 10221
rect 8095 9705 8129 9721
rect 7949 9671 8095 9705
rect 8095 9655 8129 9671
rect 16089 9705 16123 9721
rect 16123 9671 16269 9705
rect 16089 9655 16123 9671
rect 8095 9465 8129 9481
rect 7949 9431 8095 9465
rect 8095 9415 8129 9431
rect 16089 9465 16123 9481
rect 16123 9431 16269 9465
rect 16089 9415 16123 9431
rect 8095 8915 8129 8931
rect 7949 8881 8095 8915
rect 8095 8865 8129 8881
rect 16089 8915 16123 8931
rect 16123 8881 16269 8915
rect 16089 8865 16123 8881
rect 8095 8675 8129 8691
rect 7949 8641 8095 8675
rect 8095 8625 8129 8641
rect 16089 8675 16123 8691
rect 16123 8641 16269 8675
rect 16089 8625 16123 8641
rect 8095 8125 8129 8141
rect 7949 8091 8095 8125
rect 8095 8075 8129 8091
rect 16089 8125 16123 8141
rect 16123 8091 16269 8125
rect 16089 8075 16123 8091
rect 8095 7885 8129 7901
rect 7949 7851 8095 7885
rect 8095 7835 8129 7851
<< viali >>
rect 16089 14411 16123 14445
rect 8095 14171 8129 14205
rect 16089 14171 16123 14205
rect 8095 13621 8129 13655
rect 16089 13621 16123 13655
rect 8095 13381 8129 13415
rect 16089 13381 16123 13415
rect 8095 12831 8129 12865
rect 16089 12831 16123 12865
rect 8095 12591 8129 12625
rect 16089 12591 16123 12625
rect 8095 12041 8129 12075
rect 16089 12041 16123 12075
rect 8095 11801 8129 11835
rect 16089 11801 16123 11835
rect 8095 11251 8129 11285
rect 16089 11251 16123 11285
rect 8095 11011 8129 11045
rect 16089 11011 16123 11045
rect 8095 10461 8129 10495
rect 16089 10461 16123 10495
rect 8095 10221 8129 10255
rect 16089 10221 16123 10255
rect 8095 9671 8129 9705
rect 16089 9671 16123 9705
rect 8095 9431 8129 9465
rect 16089 9431 16123 9465
rect 8095 8881 8129 8915
rect 16089 8881 16123 8915
rect 8095 8641 8129 8675
rect 16089 8641 16123 8675
rect 8095 8091 8129 8125
rect 16089 8091 16123 8125
rect 8095 7851 8129 7885
<< metal1 >>
rect 9717 18358 9763 18612
rect 10711 18358 10757 18612
rect 10965 18358 11011 18612
rect 11959 18358 12005 18612
rect 12213 18358 12259 18612
rect 13207 18358 13253 18612
rect 13461 18358 13507 18612
rect 14455 18358 14501 18612
rect 14653 16202 14659 16254
rect 14711 16202 14717 16254
rect 14671 16104 14699 16202
rect 9679 15238 9707 15350
rect 10143 15238 10171 15350
rect 9679 15210 9939 15238
rect 9911 15098 9939 15210
rect 9983 15210 10171 15238
rect 10303 15238 10331 15350
rect 10767 15238 10795 15350
rect 10303 15210 10491 15238
rect 9983 15098 10011 15210
rect 10463 15098 10491 15210
rect 10535 15210 10795 15238
rect 10927 15238 10955 15350
rect 11391 15238 11419 15350
rect 10927 15210 11187 15238
rect 10535 15098 10563 15210
rect 11159 15098 11187 15210
rect 11231 15210 11419 15238
rect 11551 15238 11579 15350
rect 12015 15238 12043 15350
rect 11551 15210 11739 15238
rect 11231 15098 11259 15210
rect 11711 15098 11739 15210
rect 11783 15210 12043 15238
rect 12175 15238 12203 15350
rect 12639 15238 12667 15350
rect 12175 15210 12435 15238
rect 11783 15098 11811 15210
rect 12407 15098 12435 15210
rect 12479 15210 12667 15238
rect 12799 15238 12827 15350
rect 13263 15238 13291 15350
rect 12799 15210 12987 15238
rect 12479 15098 12507 15210
rect 12959 15098 12987 15210
rect 13031 15210 13291 15238
rect 13423 15238 13451 15350
rect 13887 15238 13915 15350
rect 13423 15210 13683 15238
rect 13031 15098 13059 15210
rect 13655 15098 13683 15210
rect 13727 15210 13915 15238
rect 14047 15238 14075 15350
rect 14511 15238 14539 15350
rect 14047 15210 14235 15238
rect 13727 15098 13755 15210
rect 14207 15098 14235 15210
rect 14279 15210 14539 15238
rect 14671 15238 14699 15350
rect 15135 15238 15163 15350
rect 14671 15210 14931 15238
rect 14279 15098 14307 15210
rect 14903 15098 14931 15210
rect 14975 15210 15163 15238
rect 14975 15098 15003 15210
rect 16074 14402 16080 14454
rect 16132 14402 16138 14454
rect 8080 14162 8086 14214
rect 8138 14162 8144 14214
rect 16074 14162 16080 14214
rect 16132 14162 16138 14214
rect 8080 13612 8086 13664
rect 8138 13612 8144 13664
rect 16074 13612 16080 13664
rect 16132 13612 16138 13664
rect 8080 13372 8086 13424
rect 8138 13372 8144 13424
rect 16074 13372 16080 13424
rect 16132 13372 16138 13424
rect 8080 12822 8086 12874
rect 8138 12822 8144 12874
rect 16074 12822 16080 12874
rect 16132 12822 16138 12874
rect 8080 12582 8086 12634
rect 8138 12582 8144 12634
rect 16074 12582 16080 12634
rect 16132 12582 16138 12634
rect 8080 12032 8086 12084
rect 8138 12032 8144 12084
rect 16074 12032 16080 12084
rect 16132 12032 16138 12084
rect 19 7988 47 11938
rect 99 7988 127 11938
rect 179 7988 207 11938
rect 259 7988 287 11938
rect 8080 11792 8086 11844
rect 8138 11792 8144 11844
rect 16074 11792 16080 11844
rect 16132 11792 16138 11844
rect 8080 11242 8086 11294
rect 8138 11242 8144 11294
rect 16074 11242 16080 11294
rect 16132 11242 16138 11294
rect 8080 11002 8086 11054
rect 8138 11002 8144 11054
rect 16074 11002 16080 11054
rect 16132 11002 16138 11054
rect 8080 10452 8086 10504
rect 8138 10452 8144 10504
rect 16074 10452 16080 10504
rect 16132 10452 16138 10504
rect 8080 10212 8086 10264
rect 8138 10212 8144 10264
rect 16074 10212 16080 10264
rect 16132 10212 16138 10264
rect 8080 9662 8086 9714
rect 8138 9662 8144 9714
rect 16074 9662 16080 9714
rect 16132 9662 16138 9714
rect 8080 9422 8086 9474
rect 8138 9422 8144 9474
rect 16074 9422 16080 9474
rect 16132 9422 16138 9474
rect 8080 8872 8086 8924
rect 8138 8872 8144 8924
rect 16074 8872 16080 8924
rect 16132 8872 16138 8924
rect 8080 8632 8086 8684
rect 8138 8632 8144 8684
rect 16074 8632 16080 8684
rect 16132 8632 16138 8684
rect 8080 8082 8086 8134
rect 8138 8082 8144 8134
rect 16074 8082 16080 8134
rect 16132 8082 16138 8134
rect 23931 7988 23959 11938
rect 24011 7988 24039 11938
rect 24091 7988 24119 11938
rect 24171 7988 24199 11938
rect 8080 7842 8086 7894
rect 8138 7842 8144 7894
rect 9431 7086 9459 7198
rect 9055 7058 9459 7086
rect 9503 7086 9531 7198
rect 9695 7086 9723 7198
rect 9503 7058 9547 7086
rect 9055 6946 9083 7058
rect 9519 6946 9547 7058
rect 9679 7058 9723 7086
rect 9767 7086 9795 7198
rect 10679 7086 10707 7198
rect 9767 7058 10171 7086
rect 9679 6946 9707 7058
rect 10143 6946 10171 7058
rect 10303 7058 10707 7086
rect 10751 7086 10779 7198
rect 10943 7086 10971 7198
rect 10751 7058 10795 7086
rect 10303 6946 10331 7058
rect 10767 6946 10795 7058
rect 10927 7058 10971 7086
rect 11015 7086 11043 7198
rect 11927 7086 11955 7198
rect 11015 7058 11419 7086
rect 10927 6946 10955 7058
rect 11391 6946 11419 7058
rect 11551 7058 11955 7086
rect 11999 7086 12027 7198
rect 12191 7086 12219 7198
rect 11999 7058 12043 7086
rect 11551 6946 11579 7058
rect 12015 6946 12043 7058
rect 12175 7058 12219 7086
rect 12263 7086 12291 7198
rect 13175 7086 13203 7198
rect 12263 7058 12667 7086
rect 12175 6946 12203 7058
rect 12639 6946 12667 7058
rect 12799 7058 13203 7086
rect 13247 7086 13275 7198
rect 13439 7086 13467 7198
rect 13247 7058 13291 7086
rect 12799 6946 12827 7058
rect 13263 6946 13291 7058
rect 13423 7058 13467 7086
rect 13511 7086 13539 7198
rect 14423 7086 14451 7198
rect 13511 7058 13915 7086
rect 13423 6946 13451 7058
rect 13887 6946 13915 7058
rect 14047 7058 14451 7086
rect 14495 7086 14523 7198
rect 14495 7058 14539 7086
rect 14047 6946 14075 7058
rect 14511 6946 14539 7058
rect 9519 6094 9547 6192
rect 9501 6042 9507 6094
rect 9559 6042 9565 6094
rect 9717 3684 9763 3938
rect 10711 3684 10757 3938
rect 10965 3684 11011 3938
rect 11959 3684 12005 3938
rect 12213 3684 12259 3938
rect 13207 3684 13253 3938
rect 13461 3684 13507 3938
rect 14455 3684 14501 3938
rect 9868 1425 9928 1481
rect 10422 1425 10482 1481
rect 11116 1425 11176 1481
rect 11670 1425 11730 1481
rect 12364 1425 12424 1481
rect 12918 1425 12978 1481
rect 13612 1425 13672 1481
rect 14166 1425 14226 1481
<< via1 >>
rect 14659 16202 14711 16254
rect 16080 14445 16132 14454
rect 16080 14411 16089 14445
rect 16089 14411 16123 14445
rect 16123 14411 16132 14445
rect 16080 14402 16132 14411
rect 8086 14205 8138 14214
rect 8086 14171 8095 14205
rect 8095 14171 8129 14205
rect 8129 14171 8138 14205
rect 8086 14162 8138 14171
rect 16080 14205 16132 14214
rect 16080 14171 16089 14205
rect 16089 14171 16123 14205
rect 16123 14171 16132 14205
rect 16080 14162 16132 14171
rect 8086 13655 8138 13664
rect 8086 13621 8095 13655
rect 8095 13621 8129 13655
rect 8129 13621 8138 13655
rect 8086 13612 8138 13621
rect 16080 13655 16132 13664
rect 16080 13621 16089 13655
rect 16089 13621 16123 13655
rect 16123 13621 16132 13655
rect 16080 13612 16132 13621
rect 8086 13415 8138 13424
rect 8086 13381 8095 13415
rect 8095 13381 8129 13415
rect 8129 13381 8138 13415
rect 8086 13372 8138 13381
rect 16080 13415 16132 13424
rect 16080 13381 16089 13415
rect 16089 13381 16123 13415
rect 16123 13381 16132 13415
rect 16080 13372 16132 13381
rect 8086 12865 8138 12874
rect 8086 12831 8095 12865
rect 8095 12831 8129 12865
rect 8129 12831 8138 12865
rect 8086 12822 8138 12831
rect 16080 12865 16132 12874
rect 16080 12831 16089 12865
rect 16089 12831 16123 12865
rect 16123 12831 16132 12865
rect 16080 12822 16132 12831
rect 8086 12625 8138 12634
rect 8086 12591 8095 12625
rect 8095 12591 8129 12625
rect 8129 12591 8138 12625
rect 8086 12582 8138 12591
rect 16080 12625 16132 12634
rect 16080 12591 16089 12625
rect 16089 12591 16123 12625
rect 16123 12591 16132 12625
rect 16080 12582 16132 12591
rect 8086 12075 8138 12084
rect 8086 12041 8095 12075
rect 8095 12041 8129 12075
rect 8129 12041 8138 12075
rect 8086 12032 8138 12041
rect 16080 12075 16132 12084
rect 16080 12041 16089 12075
rect 16089 12041 16123 12075
rect 16123 12041 16132 12075
rect 16080 12032 16132 12041
rect 8086 11835 8138 11844
rect 8086 11801 8095 11835
rect 8095 11801 8129 11835
rect 8129 11801 8138 11835
rect 8086 11792 8138 11801
rect 16080 11835 16132 11844
rect 16080 11801 16089 11835
rect 16089 11801 16123 11835
rect 16123 11801 16132 11835
rect 16080 11792 16132 11801
rect 8086 11285 8138 11294
rect 8086 11251 8095 11285
rect 8095 11251 8129 11285
rect 8129 11251 8138 11285
rect 8086 11242 8138 11251
rect 16080 11285 16132 11294
rect 16080 11251 16089 11285
rect 16089 11251 16123 11285
rect 16123 11251 16132 11285
rect 16080 11242 16132 11251
rect 8086 11045 8138 11054
rect 8086 11011 8095 11045
rect 8095 11011 8129 11045
rect 8129 11011 8138 11045
rect 8086 11002 8138 11011
rect 16080 11045 16132 11054
rect 16080 11011 16089 11045
rect 16089 11011 16123 11045
rect 16123 11011 16132 11045
rect 16080 11002 16132 11011
rect 8086 10495 8138 10504
rect 8086 10461 8095 10495
rect 8095 10461 8129 10495
rect 8129 10461 8138 10495
rect 8086 10452 8138 10461
rect 16080 10495 16132 10504
rect 16080 10461 16089 10495
rect 16089 10461 16123 10495
rect 16123 10461 16132 10495
rect 16080 10452 16132 10461
rect 8086 10255 8138 10264
rect 8086 10221 8095 10255
rect 8095 10221 8129 10255
rect 8129 10221 8138 10255
rect 8086 10212 8138 10221
rect 16080 10255 16132 10264
rect 16080 10221 16089 10255
rect 16089 10221 16123 10255
rect 16123 10221 16132 10255
rect 16080 10212 16132 10221
rect 8086 9705 8138 9714
rect 8086 9671 8095 9705
rect 8095 9671 8129 9705
rect 8129 9671 8138 9705
rect 8086 9662 8138 9671
rect 16080 9705 16132 9714
rect 16080 9671 16089 9705
rect 16089 9671 16123 9705
rect 16123 9671 16132 9705
rect 16080 9662 16132 9671
rect 8086 9465 8138 9474
rect 8086 9431 8095 9465
rect 8095 9431 8129 9465
rect 8129 9431 8138 9465
rect 8086 9422 8138 9431
rect 16080 9465 16132 9474
rect 16080 9431 16089 9465
rect 16089 9431 16123 9465
rect 16123 9431 16132 9465
rect 16080 9422 16132 9431
rect 8086 8915 8138 8924
rect 8086 8881 8095 8915
rect 8095 8881 8129 8915
rect 8129 8881 8138 8915
rect 8086 8872 8138 8881
rect 16080 8915 16132 8924
rect 16080 8881 16089 8915
rect 16089 8881 16123 8915
rect 16123 8881 16132 8915
rect 16080 8872 16132 8881
rect 8086 8675 8138 8684
rect 8086 8641 8095 8675
rect 8095 8641 8129 8675
rect 8129 8641 8138 8675
rect 8086 8632 8138 8641
rect 16080 8675 16132 8684
rect 16080 8641 16089 8675
rect 16089 8641 16123 8675
rect 16123 8641 16132 8675
rect 16080 8632 16132 8641
rect 8086 8125 8138 8134
rect 8086 8091 8095 8125
rect 8095 8091 8129 8125
rect 8129 8091 8138 8125
rect 8086 8082 8138 8091
rect 16080 8125 16132 8134
rect 16080 8091 16089 8125
rect 16089 8091 16123 8125
rect 16123 8091 16132 8125
rect 16080 8082 16132 8091
rect 8086 7885 8138 7894
rect 8086 7851 8095 7885
rect 8095 7851 8129 7885
rect 8129 7851 8138 7885
rect 8086 7842 8138 7851
rect 9507 6042 9559 6094
<< metal2 >>
rect 16289 16455 16317 18696
rect 16275 16446 16331 16455
rect 16275 16381 16331 16390
rect 14657 16256 14713 16265
rect 14657 16191 14713 16200
rect 16289 15098 16317 16381
rect 16413 16116 16441 18696
rect 16399 16107 16455 16116
rect 16399 16042 16455 16051
rect 16413 15098 16441 16042
rect 18222 14593 18250 14621
rect 16080 14454 16132 14460
rect 15979 14421 16080 14449
rect 16080 14396 16132 14402
rect 8086 14214 8138 14220
rect 16080 14214 16132 14220
rect 15979 14167 16080 14195
rect 8086 14156 8138 14162
rect 16080 14156 16132 14162
rect 8098 13975 8126 14156
rect 8098 13947 8239 13975
rect 8098 13851 8239 13879
rect 8098 13670 8126 13851
rect 8086 13664 8138 13670
rect 16080 13664 16132 13670
rect 15979 13631 16080 13659
rect 8086 13606 8138 13612
rect 16080 13606 16132 13612
rect 8086 13424 8138 13430
rect 16080 13424 16132 13430
rect 15979 13377 16080 13405
rect 8086 13366 8138 13372
rect 16080 13366 16132 13372
rect 8098 13185 8126 13366
rect 8098 13157 8239 13185
rect 8098 13061 8239 13089
rect 8098 12880 8126 13061
rect 8086 12874 8138 12880
rect 16080 12874 16132 12880
rect 15979 12841 16080 12869
rect 8086 12816 8138 12822
rect 16080 12816 16132 12822
rect 8086 12634 8138 12640
rect 16080 12634 16132 12640
rect 15979 12587 16080 12615
rect 8086 12576 8138 12582
rect 16080 12576 16132 12582
rect 8098 12395 8126 12576
rect 8098 12367 8239 12395
rect 8098 12271 8239 12299
rect 8098 12090 8126 12271
rect 8086 12084 8138 12090
rect 16080 12084 16132 12090
rect 15979 12051 16080 12079
rect 8086 12026 8138 12032
rect 16080 12026 16132 12032
rect 8086 11844 8138 11850
rect 16080 11844 16132 11850
rect 15979 11797 16080 11825
rect 8086 11786 8138 11792
rect 16080 11786 16132 11792
rect 8098 11605 8126 11786
rect 8098 11577 8239 11605
rect 8098 11481 8239 11509
rect 8098 11300 8126 11481
rect 8086 11294 8138 11300
rect 16080 11294 16132 11300
rect 15979 11261 16080 11289
rect 8086 11236 8138 11242
rect 16080 11236 16132 11242
rect 8086 11054 8138 11060
rect 16080 11054 16132 11060
rect 15979 11007 16080 11035
rect 8086 10996 8138 11002
rect 16080 10996 16132 11002
rect 8098 10815 8126 10996
rect 8098 10787 8239 10815
rect 8098 10691 8239 10719
rect 8098 10510 8126 10691
rect 8086 10504 8138 10510
rect 16080 10504 16132 10510
rect 15979 10471 16080 10499
rect 8086 10446 8138 10452
rect 16080 10446 16132 10452
rect 8086 10264 8138 10270
rect 16080 10264 16132 10270
rect 15979 10217 16080 10245
rect 8086 10206 8138 10212
rect 16080 10206 16132 10212
rect 8098 10025 8126 10206
rect 8098 9997 8239 10025
rect 8098 9901 8239 9929
rect 8098 9720 8126 9901
rect 8086 9714 8138 9720
rect 16080 9714 16132 9720
rect 15979 9681 16080 9709
rect 8086 9656 8138 9662
rect 16080 9656 16132 9662
rect 8086 9474 8138 9480
rect 16080 9474 16132 9480
rect 15979 9427 16080 9455
rect 8086 9416 8138 9422
rect 16080 9416 16132 9422
rect 8098 9235 8126 9416
rect 8098 9207 8239 9235
rect 8098 9111 8239 9139
rect 8098 8930 8126 9111
rect 8086 8924 8138 8930
rect 16080 8924 16132 8930
rect 15979 8891 16080 8919
rect 8086 8866 8138 8872
rect 16080 8866 16132 8872
rect 8086 8684 8138 8690
rect 16080 8684 16132 8690
rect 15979 8637 16080 8665
rect 8086 8626 8138 8632
rect 16080 8626 16132 8632
rect 8098 8445 8126 8626
rect 8098 8417 8239 8445
rect 8098 8321 8239 8349
rect 8098 8140 8126 8321
rect 8086 8134 8138 8140
rect 16080 8134 16132 8140
rect 15979 8101 16080 8129
rect 8086 8076 8138 8082
rect 16080 8076 16132 8082
rect 8086 7894 8138 7900
rect 8086 7836 8138 7842
rect 5968 7675 5996 7703
rect 8098 7655 8126 7836
rect 8098 7627 8239 7655
rect 7619 6254 7647 7198
rect 7605 6245 7661 6254
rect 7605 6180 7661 6189
rect 7619 49 7647 6180
rect 7743 5915 7771 7198
rect 7729 5906 7785 5915
rect 7729 5841 7785 5850
rect 7743 49 7771 5841
rect 7867 604 7895 7198
rect 9505 6096 9561 6105
rect 9505 6031 9561 6040
rect 7853 595 7909 604
rect 7853 530 7909 539
rect 7867 49 7895 530
rect 9599 305 9627 333
rect 10847 305 10875 333
rect 12095 305 12123 333
rect 13343 305 13371 333
<< via2 >>
rect 16275 16390 16331 16446
rect 14657 16254 14713 16256
rect 14657 16202 14659 16254
rect 14659 16202 14711 16254
rect 14711 16202 14713 16254
rect 14657 16200 14713 16202
rect 16399 16051 16455 16107
rect 7605 6189 7661 6245
rect 7729 5850 7785 5906
rect 9505 6094 9561 6096
rect 9505 6042 9507 6094
rect 9507 6042 9559 6094
rect 9559 6042 9561 6094
rect 9505 6040 9561 6042
rect 7853 539 7909 595
<< metal3 >>
rect 9945 18455 10043 18553
rect 10431 18455 10529 18553
rect 11193 18455 11291 18553
rect 11679 18455 11777 18553
rect 12441 18455 12539 18553
rect 12927 18455 13025 18553
rect 13689 18455 13787 18553
rect 14175 18455 14273 18553
rect 9945 18133 10043 18231
rect 10431 18133 10529 18231
rect 11193 18133 11291 18231
rect 11679 18133 11777 18231
rect 12441 18133 12539 18231
rect 12927 18133 13025 18231
rect 13689 18133 13787 18231
rect 14175 18133 14273 18231
rect 9933 17295 10031 17393
rect 10443 17295 10541 17393
rect 11181 17295 11279 17393
rect 11691 17295 11789 17393
rect 12429 17295 12527 17393
rect 12939 17295 13037 17393
rect 13677 17295 13775 17393
rect 14187 17295 14285 17393
rect 10015 16521 10113 16619
rect 10361 16521 10459 16619
rect 11263 16521 11361 16619
rect 11609 16521 11707 16619
rect 12511 16521 12609 16619
rect 12857 16521 12955 16619
rect 13759 16521 13857 16619
rect 14105 16521 14203 16619
rect 16270 16448 16336 16451
rect 11422 16446 16336 16448
rect 11422 16390 16275 16446
rect 16331 16390 16336 16446
rect 11422 16388 16336 16390
rect 16270 16385 16336 16388
rect 14652 16258 14718 16261
rect 14652 16256 24302 16258
rect 14652 16200 14657 16256
rect 14713 16200 24302 16256
rect 14652 16198 24302 16200
rect 14652 16195 14718 16198
rect 16394 16109 16460 16112
rect 11734 16107 16460 16109
rect 11734 16051 16399 16107
rect 16455 16051 16460 16107
rect 11734 16049 16460 16051
rect 16394 16046 16460 16049
rect 9757 15411 9855 15509
rect 10619 15411 10717 15509
rect 11005 15411 11103 15509
rect 11867 15411 11965 15509
rect 12253 15411 12351 15509
rect 13115 15411 13213 15509
rect 13501 15411 13599 15509
rect 14363 15411 14461 15509
rect 14749 15411 14847 15509
rect 9252 14820 9350 14918
rect 9876 14820 9974 14918
rect 10500 14820 10598 14918
rect 11124 14820 11222 14918
rect 11748 14820 11846 14918
rect 12372 14820 12470 14918
rect 12996 14820 13094 14918
rect 13620 14820 13718 14918
rect 14244 14820 14342 14918
rect 14868 14820 14966 14918
rect 8190 14606 8288 14704
rect 15930 14606 16028 14704
rect 16556 14456 16654 14554
rect 17595 14444 17693 14542
rect 18427 14450 18525 14548
rect 8556 14259 8654 14357
rect 15564 14259 15662 14357
rect 8556 14022 8654 14120
rect 15564 14022 15662 14120
rect 4468 13871 4566 13969
rect 4893 13871 4991 13969
rect 5272 13864 5370 13962
rect 5668 13864 5766 13962
rect 18452 13864 18550 13962
rect 18848 13864 18946 13962
rect 19227 13871 19325 13969
rect 19652 13871 19750 13969
rect 8556 13706 8654 13804
rect 15564 13706 15662 13804
rect 4468 13499 4566 13597
rect 4893 13501 4991 13599
rect 5272 13469 5370 13567
rect 5668 13469 5766 13567
rect 8556 13469 8654 13567
rect 15564 13469 15662 13567
rect 18452 13469 18550 13567
rect 18848 13469 18946 13567
rect 19227 13501 19325 13599
rect 19652 13499 19750 13597
rect 8556 13232 8654 13330
rect 15564 13232 15662 13330
rect 4468 13081 4566 13179
rect 4893 13081 4991 13179
rect 5272 13074 5370 13172
rect 5668 13074 5766 13172
rect 18452 13074 18550 13172
rect 18848 13074 18946 13172
rect 19227 13081 19325 13179
rect 19652 13081 19750 13179
rect 8556 12916 8654 13014
rect 15564 12916 15662 13014
rect 4468 12709 4566 12807
rect 4893 12711 4991 12809
rect 5272 12679 5370 12777
rect 5668 12679 5766 12777
rect 8556 12679 8654 12777
rect 15564 12679 15662 12777
rect 18452 12679 18550 12777
rect 18848 12679 18946 12777
rect 19227 12711 19325 12809
rect 19652 12709 19750 12807
rect 8556 12442 8654 12540
rect 15564 12442 15662 12540
rect 4468 12291 4566 12389
rect 4893 12291 4991 12389
rect 5272 12284 5370 12382
rect 5668 12284 5766 12382
rect 18452 12284 18550 12382
rect 18848 12284 18946 12382
rect 19227 12291 19325 12389
rect 19652 12291 19750 12389
rect 8556 12126 8654 12224
rect 15564 12126 15662 12224
rect 4468 11919 4566 12017
rect 4893 11921 4991 12019
rect 5272 11889 5370 11987
rect 5668 11889 5766 11987
rect 8556 11889 8654 11987
rect 15564 11889 15662 11987
rect 18452 11889 18550 11987
rect 18848 11889 18946 11987
rect 19227 11921 19325 12019
rect 19652 11919 19750 12017
rect 8556 11652 8654 11750
rect 15564 11652 15662 11750
rect 2130 11501 2228 11599
rect 2555 11501 2653 11599
rect 2934 11494 3032 11592
rect 3330 11494 3428 11592
rect 4468 11501 4566 11599
rect 4893 11501 4991 11599
rect 5272 11494 5370 11592
rect 5668 11494 5766 11592
rect 18452 11494 18550 11592
rect 18848 11494 18946 11592
rect 19227 11501 19325 11599
rect 19652 11501 19750 11599
rect 20790 11494 20888 11592
rect 21186 11494 21284 11592
rect 21565 11501 21663 11599
rect 21990 11501 22088 11599
rect 8556 11336 8654 11434
rect 15564 11336 15662 11434
rect 4468 11129 4566 11227
rect 4893 11131 4991 11229
rect 5272 11099 5370 11197
rect 5668 11099 5766 11197
rect 6100 11084 6198 11182
rect 6525 11083 6623 11181
rect 6942 11099 7040 11197
rect 7564 11099 7662 11197
rect 8556 11099 8654 11197
rect 15564 11099 15662 11197
rect 16556 11099 16654 11197
rect 17178 11099 17276 11197
rect 17595 11083 17693 11181
rect 18020 11084 18118 11182
rect 18452 11099 18550 11197
rect 18848 11099 18946 11197
rect 19227 11131 19325 11229
rect 19652 11129 19750 11227
rect 8556 10862 8654 10960
rect 15564 10862 15662 10960
rect 836 10704 934 10802
rect 1232 10704 1330 10802
rect 2130 10711 2228 10809
rect 2555 10711 2653 10809
rect 2934 10704 3032 10802
rect 3330 10704 3428 10802
rect 4468 10711 4566 10809
rect 4893 10711 4991 10809
rect 5272 10704 5370 10802
rect 5668 10704 5766 10802
rect 18452 10704 18550 10802
rect 18848 10704 18946 10802
rect 19227 10711 19325 10809
rect 19652 10711 19750 10809
rect 20790 10704 20888 10802
rect 21186 10704 21284 10802
rect 21565 10711 21663 10809
rect 21990 10711 22088 10809
rect 22888 10704 22986 10802
rect 23284 10704 23382 10802
rect 8556 10546 8654 10644
rect 15564 10546 15662 10644
rect 4468 10339 4566 10437
rect 4893 10341 4991 10439
rect 5272 10309 5370 10407
rect 5668 10309 5766 10407
rect 8556 10309 8654 10407
rect 15564 10309 15662 10407
rect 18452 10309 18550 10407
rect 18848 10309 18946 10407
rect 19227 10341 19325 10439
rect 19652 10339 19750 10437
rect 8556 10072 8654 10170
rect 15564 10072 15662 10170
rect 4468 9921 4566 10019
rect 4893 9921 4991 10019
rect 5272 9914 5370 10012
rect 5668 9914 5766 10012
rect 18452 9914 18550 10012
rect 18848 9914 18946 10012
rect 19227 9921 19325 10019
rect 19652 9921 19750 10019
rect 8556 9756 8654 9854
rect 15564 9756 15662 9854
rect 4468 9549 4566 9647
rect 4893 9551 4991 9649
rect 5272 9519 5370 9617
rect 5668 9519 5766 9617
rect 8556 9519 8654 9617
rect 15564 9519 15662 9617
rect 18452 9519 18550 9617
rect 18848 9519 18946 9617
rect 19227 9551 19325 9649
rect 19652 9549 19750 9647
rect 8556 9282 8654 9380
rect 15564 9282 15662 9380
rect 2130 9131 2228 9229
rect 2555 9131 2653 9229
rect 2934 9124 3032 9222
rect 3330 9124 3428 9222
rect 4468 9131 4566 9229
rect 4893 9131 4991 9229
rect 5272 9124 5370 9222
rect 5668 9124 5766 9222
rect 18452 9124 18550 9222
rect 18848 9124 18946 9222
rect 19227 9131 19325 9229
rect 19652 9131 19750 9229
rect 20790 9124 20888 9222
rect 21186 9124 21284 9222
rect 21565 9131 21663 9229
rect 21990 9131 22088 9229
rect 8556 8966 8654 9064
rect 15564 8966 15662 9064
rect 4468 8759 4566 8857
rect 4893 8761 4991 8859
rect 5272 8729 5370 8827
rect 5668 8729 5766 8827
rect 8556 8729 8654 8827
rect 15564 8729 15662 8827
rect 18452 8729 18550 8827
rect 18848 8729 18946 8827
rect 19227 8761 19325 8859
rect 19652 8759 19750 8857
rect 8556 8492 8654 8590
rect 15564 8492 15662 8590
rect 836 8334 934 8432
rect 1232 8334 1330 8432
rect 2130 8341 2228 8439
rect 2555 8341 2653 8439
rect 2934 8334 3032 8432
rect 3330 8334 3428 8432
rect 4468 8341 4566 8439
rect 4893 8341 4991 8439
rect 5272 8334 5370 8432
rect 5668 8334 5766 8432
rect 18452 8334 18550 8432
rect 18848 8334 18946 8432
rect 19227 8341 19325 8439
rect 19652 8341 19750 8439
rect 20790 8334 20888 8432
rect 21186 8334 21284 8432
rect 21565 8341 21663 8439
rect 21990 8341 22088 8439
rect 22888 8334 22986 8432
rect 23284 8334 23382 8432
rect 8556 8176 8654 8274
rect 15564 8176 15662 8274
rect 8556 7939 8654 8037
rect 15564 7939 15662 8037
rect 5693 7748 5791 7846
rect 6525 7754 6623 7852
rect 7564 7742 7662 7840
rect 8190 7812 8288 7910
rect 15930 7812 16028 7910
rect 9252 7378 9350 7476
rect 9876 7378 9974 7476
rect 10500 7378 10598 7476
rect 11124 7378 11222 7476
rect 11748 7378 11846 7476
rect 12372 7378 12470 7476
rect 12996 7378 13094 7476
rect 13620 7378 13718 7476
rect 14244 7378 14342 7476
rect 14868 7378 14966 7476
rect 9371 6787 9469 6885
rect 9757 6787 9855 6885
rect 10619 6787 10717 6885
rect 11005 6787 11103 6885
rect 11867 6787 11965 6885
rect 12253 6787 12351 6885
rect 13115 6787 13213 6885
rect 13501 6787 13599 6885
rect 14363 6787 14461 6885
rect 7600 6247 7666 6250
rect 7600 6245 11422 6247
rect 7600 6189 7605 6245
rect 7661 6189 11422 6245
rect 7600 6187 11422 6189
rect 7600 6184 7666 6187
rect 9500 6098 9566 6101
rect 0 6096 9566 6098
rect 0 6040 9505 6096
rect 9561 6040 9566 6096
rect 0 6038 9566 6040
rect 9500 6035 9566 6038
rect 7724 5908 7790 5911
rect 7724 5906 11422 5908
rect 7724 5850 7729 5906
rect 7785 5850 11422 5906
rect 7724 5848 11422 5850
rect 7724 5845 7790 5848
rect 10015 5677 10113 5775
rect 10361 5677 10459 5775
rect 11263 5677 11361 5775
rect 11609 5677 11707 5775
rect 12511 5677 12609 5775
rect 12857 5677 12955 5775
rect 13759 5677 13857 5775
rect 14105 5677 14203 5775
rect 9933 4903 10031 5001
rect 10443 4903 10541 5001
rect 11181 4903 11279 5001
rect 11691 4903 11789 5001
rect 12429 4903 12527 5001
rect 12939 4903 13037 5001
rect 13677 4903 13775 5001
rect 14187 4903 14285 5001
rect 9945 4065 10043 4163
rect 10431 4065 10529 4163
rect 11193 4065 11291 4163
rect 11679 4065 11777 4163
rect 12441 4065 12539 4163
rect 12927 4065 13025 4163
rect 13689 4065 13787 4163
rect 14175 4065 14273 4163
rect 9945 3743 10043 3841
rect 10431 3743 10529 3841
rect 11193 3743 11291 3841
rect 11679 3743 11777 3841
rect 12441 3743 12539 3841
rect 12927 3743 13025 3841
rect 13689 3743 13787 3841
rect 14175 3743 14273 3841
rect 9831 2950 9929 3048
rect 10421 2950 10519 3048
rect 11079 2950 11177 3048
rect 11669 2950 11767 3048
rect 12327 2950 12425 3048
rect 12917 2950 13015 3048
rect 13575 2950 13673 3048
rect 14165 2950 14263 3048
rect 9820 2513 9918 2611
rect 10432 2513 10530 2611
rect 11068 2513 11166 2611
rect 11680 2513 11778 2611
rect 12316 2513 12414 2611
rect 12928 2513 13026 2611
rect 13564 2513 13662 2611
rect 14176 2513 14274 2611
rect 9941 2181 10039 2279
rect 10311 2181 10409 2279
rect 11189 2181 11287 2279
rect 11559 2181 11657 2279
rect 12437 2181 12535 2279
rect 12807 2181 12905 2279
rect 13685 2181 13783 2279
rect 14055 2181 14153 2279
rect 9826 1979 9924 2077
rect 10426 1979 10524 2077
rect 11074 1979 11172 2077
rect 11674 1979 11772 2077
rect 12322 1979 12420 2077
rect 12922 1979 13020 2077
rect 13570 1979 13668 2077
rect 14170 1979 14268 2077
rect 9840 1563 9938 1661
rect 10412 1563 10510 1661
rect 11088 1563 11186 1661
rect 11660 1563 11758 1661
rect 12336 1563 12434 1661
rect 12908 1563 13006 1661
rect 13584 1563 13682 1661
rect 14156 1563 14254 1661
rect 8190 1120 8288 1218
rect 14556 1120 14654 1218
rect 7848 597 7914 600
rect 7848 595 11422 597
rect 7848 539 7853 595
rect 7909 539 11422 595
rect 7848 537 11422 539
rect 7848 534 7914 537
rect 8190 0 8288 98
rect 14556 0 14654 98
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 16270 0 1 16381
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 16394 0 1 16042
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 16074 0 1 14396
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 16077 0 1 14395
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 16074 0 1 14156
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 16077 0 1 14155
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 16074 0 1 13606
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 16077 0 1 13605
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 16074 0 1 13366
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 16077 0 1 13365
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 16074 0 1 12816
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 16077 0 1 12815
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 16074 0 1 12576
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 16077 0 1 12575
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 16074 0 1 12026
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 16077 0 1 12025
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 16074 0 1 11786
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 16077 0 1 11785
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 16074 0 1 11236
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 16077 0 1 11235
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 16074 0 1 10996
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 16077 0 1 10995
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 16074 0 1 10446
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 16077 0 1 10445
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 16074 0 1 10206
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 16077 0 1 10205
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 16074 0 1 9656
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1634918361
transform 1 0 16077 0 1 9655
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 16074 0 1 9416
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1634918361
transform 1 0 16077 0 1 9415
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 16074 0 1 8866
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1634918361
transform 1 0 16077 0 1 8865
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 16074 0 1 8626
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1634918361
transform 1 0 16077 0 1 8625
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1634918361
transform 1 0 16074 0 1 8076
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1634918361
transform 1 0 16077 0 1 8075
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 14652 0 1 16191
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1634918361
transform 1 0 14653 0 1 16196
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 7724 0 1 5841
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 7848 0 1 530
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 7600 0 1 6180
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1634918361
transform 1 0 8080 0 1 7836
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1634918361
transform 1 0 8083 0 1 7835
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1634918361
transform 1 0 8080 0 1 14156
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1634918361
transform 1 0 8083 0 1 14155
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1634918361
transform 1 0 8080 0 1 13606
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1634918361
transform 1 0 8083 0 1 13605
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1634918361
transform 1 0 8080 0 1 13366
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1634918361
transform 1 0 8083 0 1 13365
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1634918361
transform 1 0 8080 0 1 12816
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1634918361
transform 1 0 8083 0 1 12815
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1634918361
transform 1 0 8080 0 1 12576
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1634918361
transform 1 0 8083 0 1 12575
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1634918361
transform 1 0 8080 0 1 12026
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1634918361
transform 1 0 8083 0 1 12025
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1634918361
transform 1 0 8080 0 1 11786
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1634918361
transform 1 0 8083 0 1 11785
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1634918361
transform 1 0 8080 0 1 11236
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1634918361
transform 1 0 8083 0 1 11235
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1634918361
transform 1 0 8080 0 1 10996
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1634918361
transform 1 0 8083 0 1 10995
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1634918361
transform 1 0 8080 0 1 10446
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1634918361
transform 1 0 8083 0 1 10445
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1634918361
transform 1 0 8080 0 1 10206
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1634918361
transform 1 0 8083 0 1 10205
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1634918361
transform 1 0 8080 0 1 9656
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1634918361
transform 1 0 8083 0 1 9655
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1634918361
transform 1 0 8080 0 1 9416
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1634918361
transform 1 0 8083 0 1 9415
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1634918361
transform 1 0 8080 0 1 8866
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1634918361
transform 1 0 8083 0 1 8865
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1634918361
transform 1 0 8080 0 1 8626
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1634918361
transform 1 0 8083 0 1 8625
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1634918361
transform 1 0 8080 0 1 8076
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1634918361
transform 1 0 8083 0 1 8075
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 9500 0 1 6031
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1634918361
transform 1 0 9501 0 1 6036
box 0 0 1 1
use port_address_0  port_address_0_0
timestamp 1634918361
transform -1 0 24218 0 1 7988
box 0 -56 7967 6810
use port_address  port_address_0
timestamp 1634918361
transform 1 0 0 0 1 7988
box 0 -490 7967 6376
use port_data_0  port_data_0_0
timestamp 1634918361
transform 1 0 8239 0 1 15098
box 0 238 6990 3514
use port_data  port_data_0
timestamp 1634918361
transform 1 0 8239 0 -1 7198
box -49 238 6907 7198
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1634918361
transform 1 0 8239 0 1 7198
box -49 0 7789 7900
<< labels >>
rlabel metal2 s 7619 49 7647 7198 4 p_en_bar0
port 1 nsew
rlabel metal2 s 7743 49 7771 7198 4 s_en0
port 2 nsew
rlabel metal2 s 7867 49 7895 7198 4 w_en0
port 3 nsew
rlabel metal2 s 5968 7675 5996 7703 4 wl_en0
port 4 nsew
rlabel metal2 s 16289 15098 16317 18696 4 s_en1
port 5 nsew
rlabel metal2 s 16413 15098 16441 18696 4 p_en_bar1
port 6 nsew
rlabel metal2 s 18222 14593 18250 14621 4 wl_en1
port 7 nsew
rlabel metal1 s 9868 1425 9928 1481 4 din0_0
port 8 nsew
rlabel metal1 s 10422 1425 10482 1481 4 din0_1
port 9 nsew
rlabel metal1 s 11116 1425 11176 1481 4 din0_2
port 10 nsew
rlabel metal1 s 11670 1425 11730 1481 4 din0_3
port 11 nsew
rlabel metal1 s 12364 1425 12424 1481 4 din0_4
port 12 nsew
rlabel metal1 s 12918 1425 12978 1481 4 din0_5
port 13 nsew
rlabel metal1 s 13612 1425 13672 1481 4 din0_6
port 14 nsew
rlabel metal1 s 14166 1425 14226 1481 4 din0_7
port 15 nsew
rlabel metal2 s 9599 305 9627 333 4 bank_wmask0_0
port 16 nsew
rlabel metal2 s 10847 305 10875 333 4 bank_wmask0_1
port 17 nsew
rlabel metal2 s 12095 305 12123 333 4 bank_wmask0_2
port 18 nsew
rlabel metal2 s 13343 305 13371 333 4 bank_wmask0_3
port 19 nsew
rlabel metal1 s 9717 3684 9763 3938 4 dout0_0
port 20 nsew
rlabel metal1 s 10711 3684 10757 3938 4 dout0_1
port 21 nsew
rlabel metal1 s 10965 3684 11011 3938 4 dout0_2
port 22 nsew
rlabel metal1 s 11959 3684 12005 3938 4 dout0_3
port 23 nsew
rlabel metal1 s 12213 3684 12259 3938 4 dout0_4
port 24 nsew
rlabel metal1 s 13207 3684 13253 3938 4 dout0_5
port 25 nsew
rlabel metal1 s 13461 3684 13507 3938 4 dout0_6
port 26 nsew
rlabel metal1 s 14455 3684 14501 3938 4 dout0_7
port 27 nsew
rlabel metal3 s 0 6038 9533 6098 4 rbl_bl_0_0
port 28 nsew
rlabel metal1 s 19 7988 47 11938 4 addr0_0
port 29 nsew
rlabel metal1 s 99 7988 127 11938 4 addr0_1
port 30 nsew
rlabel metal1 s 179 7988 207 11938 4 addr0_2
port 31 nsew
rlabel metal1 s 259 7988 287 11938 4 addr0_3
port 32 nsew
rlabel metal1 s 9717 18358 9763 18612 4 dout1_0
port 33 nsew
rlabel metal1 s 10711 18358 10757 18612 4 dout1_1
port 34 nsew
rlabel metal1 s 10965 18358 11011 18612 4 dout1_2
port 35 nsew
rlabel metal1 s 11959 18358 12005 18612 4 dout1_3
port 36 nsew
rlabel metal1 s 12213 18358 12259 18612 4 dout1_4
port 37 nsew
rlabel metal1 s 13207 18358 13253 18612 4 dout1_5
port 38 nsew
rlabel metal1 s 13461 18358 13507 18612 4 dout1_6
port 39 nsew
rlabel metal1 s 14455 18358 14501 18612 4 dout1_7
port 40 nsew
rlabel metal3 s 14685 16198 24302 16258 4 rbl_bl_1_1
port 41 nsew
rlabel metal1 s 24171 7988 24199 11938 4 addr1_0
port 42 nsew
rlabel metal1 s 24091 7988 24119 11938 4 addr1_1
port 43 nsew
rlabel metal1 s 24011 7988 24039 11938 4 addr1_2
port 44 nsew
rlabel metal1 s 23931 7988 23959 11938 4 addr1_3
port 45 nsew
rlabel metal3 s 19227 9131 19325 9229 4 vdd
port 46 nsew
rlabel metal3 s 4893 8761 4991 8859 4 vdd
port 46 nsew
rlabel metal3 s 4893 12711 4991 12809 4 vdd
port 46 nsew
rlabel metal3 s 9252 7378 9350 7476 4 vdd
port 46 nsew
rlabel metal3 s 17595 11083 17693 11181 4 vdd
port 46 nsew
rlabel metal3 s 12927 18133 13025 18231 4 vdd
port 46 nsew
rlabel metal3 s 4893 10341 4991 10439 4 vdd
port 46 nsew
rlabel metal3 s 9840 1563 9938 1661 4 vdd
port 46 nsew
rlabel metal3 s 5668 11889 5766 11987 4 vdd
port 46 nsew
rlabel metal3 s 14187 17295 14285 17393 4 vdd
port 46 nsew
rlabel metal3 s 18452 12284 18550 12382 4 vdd
port 46 nsew
rlabel metal3 s 21565 8341 21663 8439 4 vdd
port 46 nsew
rlabel metal3 s 14176 2513 14274 2611 4 vdd
port 46 nsew
rlabel metal3 s 3330 11494 3428 11592 4 vdd
port 46 nsew
rlabel metal3 s 9876 7378 9974 7476 4 vdd
port 46 nsew
rlabel metal3 s 10432 2513 10530 2611 4 vdd
port 46 nsew
rlabel metal3 s 11691 4903 11789 5001 4 vdd
port 46 nsew
rlabel metal3 s 11181 17295 11279 17393 4 vdd
port 46 nsew
rlabel metal3 s 10619 15411 10717 15509 4 vdd
port 46 nsew
rlabel metal3 s 4893 9131 4991 9229 4 vdd
port 46 nsew
rlabel metal3 s 12908 1563 13006 1661 4 vdd
port 46 nsew
rlabel metal3 s 5668 9124 5766 9222 4 vdd
port 46 nsew
rlabel metal3 s 18452 12679 18550 12777 4 vdd
port 46 nsew
rlabel metal3 s 4893 10711 4991 10809 4 vdd
port 46 nsew
rlabel metal3 s 11679 4065 11777 4163 4 vdd
port 46 nsew
rlabel metal3 s 19227 8761 19325 8859 4 vdd
port 46 nsew
rlabel metal3 s 11660 1563 11758 1661 4 vdd
port 46 nsew
rlabel metal3 s 18452 11099 18550 11197 4 vdd
port 46 nsew
rlabel metal3 s 18452 9124 18550 9222 4 vdd
port 46 nsew
rlabel metal3 s 3330 8334 3428 8432 4 vdd
port 46 nsew
rlabel metal3 s 4893 9551 4991 9649 4 vdd
port 46 nsew
rlabel metal3 s 14556 1120 14654 1218 4 vdd
port 46 nsew
rlabel metal3 s 9820 2513 9918 2611 4 vdd
port 46 nsew
rlabel metal3 s 4893 8341 4991 8439 4 vdd
port 46 nsew
rlabel metal3 s 21565 11501 21663 11599 4 vdd
port 46 nsew
rlabel metal3 s 19227 13501 19325 13599 4 vdd
port 46 nsew
rlabel metal3 s 6525 11083 6623 11181 4 vdd
port 46 nsew
rlabel metal3 s 14749 15411 14847 15509 4 vdd
port 46 nsew
rlabel metal3 s 12372 7378 12470 7476 4 vdd
port 46 nsew
rlabel metal3 s 5693 7748 5791 7846 4 vdd
port 46 nsew
rlabel metal3 s 13677 4903 13775 5001 4 vdd
port 46 nsew
rlabel metal3 s 12441 18133 12539 18231 4 vdd
port 46 nsew
rlabel metal3 s 13115 15411 13213 15509 4 vdd
port 46 nsew
rlabel metal3 s 18452 13864 18550 13962 4 vdd
port 46 nsew
rlabel metal3 s 13689 18133 13787 18231 4 vdd
port 46 nsew
rlabel metal3 s 4893 11501 4991 11599 4 vdd
port 46 nsew
rlabel metal3 s 16556 14456 16654 14554 4 vdd
port 46 nsew
rlabel metal3 s 12372 14820 12470 14918 4 vdd
port 46 nsew
rlabel metal3 s 11193 4065 11291 4163 4 vdd
port 46 nsew
rlabel metal3 s 16556 11099 16654 11197 4 vdd
port 46 nsew
rlabel metal3 s 18452 13469 18550 13567 4 vdd
port 46 nsew
rlabel metal3 s 11867 6787 11965 6885 4 vdd
port 46 nsew
rlabel metal3 s 19227 13081 19325 13179 4 vdd
port 46 nsew
rlabel metal3 s 21565 10711 21663 10809 4 vdd
port 46 nsew
rlabel metal3 s 5668 11494 5766 11592 4 vdd
port 46 nsew
rlabel metal3 s 13689 4065 13787 4163 4 vdd
port 46 nsew
rlabel metal3 s 20790 11494 20888 11592 4 vdd
port 46 nsew
rlabel metal3 s 18452 11494 18550 11592 4 vdd
port 46 nsew
rlabel metal3 s 10500 14820 10598 14918 4 vdd
port 46 nsew
rlabel metal3 s 5668 9519 5766 9617 4 vdd
port 46 nsew
rlabel metal3 s 11691 17295 11789 17393 4 vdd
port 46 nsew
rlabel metal3 s 17595 14444 17693 14542 4 vdd
port 46 nsew
rlabel metal3 s 11679 18133 11777 18231 4 vdd
port 46 nsew
rlabel metal3 s 4893 12291 4991 12389 4 vdd
port 46 nsew
rlabel metal3 s 12429 4903 12527 5001 4 vdd
port 46 nsew
rlabel metal3 s 9876 14820 9974 14918 4 vdd
port 46 nsew
rlabel metal3 s 12939 17295 13037 17393 4 vdd
port 46 nsew
rlabel metal3 s 5668 10309 5766 10407 4 vdd
port 46 nsew
rlabel metal3 s 12996 14820 13094 14918 4 vdd
port 46 nsew
rlabel metal3 s 14244 7378 14342 7476 4 vdd
port 46 nsew
rlabel metal3 s 14244 14820 14342 14918 4 vdd
port 46 nsew
rlabel metal3 s 14363 6787 14461 6885 4 vdd
port 46 nsew
rlabel metal3 s 14156 1563 14254 1661 4 vdd
port 46 nsew
rlabel metal3 s 12928 2513 13026 2611 4 vdd
port 46 nsew
rlabel metal3 s 4893 11131 4991 11229 4 vdd
port 46 nsew
rlabel metal3 s 20790 8334 20888 8432 4 vdd
port 46 nsew
rlabel metal3 s 5668 8729 5766 8827 4 vdd
port 46 nsew
rlabel metal3 s 10500 7378 10598 7476 4 vdd
port 46 nsew
rlabel metal3 s 18452 8334 18550 8432 4 vdd
port 46 nsew
rlabel metal3 s 9933 17295 10031 17393 4 vdd
port 46 nsew
rlabel metal3 s 10443 4903 10541 5001 4 vdd
port 46 nsew
rlabel metal3 s 11068 2513 11166 2611 4 vdd
port 46 nsew
rlabel metal3 s 4893 13081 4991 13179 4 vdd
port 46 nsew
rlabel metal3 s 19227 11501 19325 11599 4 vdd
port 46 nsew
rlabel metal3 s 14187 4903 14285 5001 4 vdd
port 46 nsew
rlabel metal3 s 11867 15411 11965 15509 4 vdd
port 46 nsew
rlabel metal3 s 9252 14820 9350 14918 4 vdd
port 46 nsew
rlabel metal3 s 18452 10704 18550 10802 4 vdd
port 46 nsew
rlabel metal3 s 11005 6787 11103 6885 4 vdd
port 46 nsew
rlabel metal3 s 10619 6787 10717 6885 4 vdd
port 46 nsew
rlabel metal3 s 4893 9921 4991 10019 4 vdd
port 46 nsew
rlabel metal3 s 13501 6787 13599 6885 4 vdd
port 46 nsew
rlabel metal3 s 9945 18133 10043 18231 4 vdd
port 46 nsew
rlabel metal3 s 14363 15411 14461 15509 4 vdd
port 46 nsew
rlabel metal3 s 5668 13864 5766 13962 4 vdd
port 46 nsew
rlabel metal3 s 2555 10711 2653 10809 4 vdd
port 46 nsew
rlabel metal3 s 18452 9519 18550 9617 4 vdd
port 46 nsew
rlabel metal3 s 9371 6787 9469 6885 4 vdd
port 46 nsew
rlabel metal3 s 18452 10309 18550 10407 4 vdd
port 46 nsew
rlabel metal3 s 7564 11099 7662 11197 4 vdd
port 46 nsew
rlabel metal3 s 5668 13074 5766 13172 4 vdd
port 46 nsew
rlabel metal3 s 13620 14820 13718 14918 4 vdd
port 46 nsew
rlabel metal3 s 12336 1563 12434 1661 4 vdd
port 46 nsew
rlabel metal3 s 11124 7378 11222 7476 4 vdd
port 46 nsew
rlabel metal3 s 3330 9124 3428 9222 4 vdd
port 46 nsew
rlabel metal3 s 10431 4065 10529 4163 4 vdd
port 46 nsew
rlabel metal3 s 11181 4903 11279 5001 4 vdd
port 46 nsew
rlabel metal3 s 2555 8341 2653 8439 4 vdd
port 46 nsew
rlabel metal3 s 19227 12711 19325 12809 4 vdd
port 46 nsew
rlabel metal3 s 11088 1563 11186 1661 4 vdd
port 46 nsew
rlabel metal3 s 14868 7378 14966 7476 4 vdd
port 46 nsew
rlabel metal3 s 8190 1120 8288 1218 4 vdd
port 46 nsew
rlabel metal3 s 10443 17295 10541 17393 4 vdd
port 46 nsew
rlabel metal3 s 19227 9551 19325 9649 4 vdd
port 46 nsew
rlabel metal3 s 12429 17295 12527 17393 4 vdd
port 46 nsew
rlabel metal3 s 14868 14820 14966 14918 4 vdd
port 46 nsew
rlabel metal3 s 19227 8341 19325 8439 4 vdd
port 46 nsew
rlabel metal3 s 2555 11501 2653 11599 4 vdd
port 46 nsew
rlabel metal3 s 18452 11889 18550 11987 4 vdd
port 46 nsew
rlabel metal3 s 14175 4065 14273 4163 4 vdd
port 46 nsew
rlabel metal3 s 10412 1563 10510 1661 4 vdd
port 46 nsew
rlabel metal3 s 1232 8334 1330 8432 4 vdd
port 46 nsew
rlabel metal3 s 12996 7378 13094 7476 4 vdd
port 46 nsew
rlabel metal3 s 19227 10711 19325 10809 4 vdd
port 46 nsew
rlabel metal3 s 9945 4065 10043 4163 4 vdd
port 46 nsew
rlabel metal3 s 22888 10704 22986 10802 4 vdd
port 46 nsew
rlabel metal3 s 18452 13074 18550 13172 4 vdd
port 46 nsew
rlabel metal3 s 5668 9914 5766 10012 4 vdd
port 46 nsew
rlabel metal3 s 13564 2513 13662 2611 4 vdd
port 46 nsew
rlabel metal3 s 9757 6787 9855 6885 4 vdd
port 46 nsew
rlabel metal3 s 4893 13501 4991 13599 4 vdd
port 46 nsew
rlabel metal3 s 13115 6787 13213 6885 4 vdd
port 46 nsew
rlabel metal3 s 5668 13469 5766 13567 4 vdd
port 46 nsew
rlabel metal3 s 10431 18133 10529 18231 4 vdd
port 46 nsew
rlabel metal3 s 11680 2513 11778 2611 4 vdd
port 46 nsew
rlabel metal3 s 18452 9914 18550 10012 4 vdd
port 46 nsew
rlabel metal3 s 11005 15411 11103 15509 4 vdd
port 46 nsew
rlabel metal3 s 20790 9124 20888 9222 4 vdd
port 46 nsew
rlabel metal3 s 4893 11921 4991 12019 4 vdd
port 46 nsew
rlabel metal3 s 11748 14820 11846 14918 4 vdd
port 46 nsew
rlabel metal3 s 3330 10704 3428 10802 4 vdd
port 46 nsew
rlabel metal3 s 19227 10341 19325 10439 4 vdd
port 46 nsew
rlabel metal3 s 12316 2513 12414 2611 4 vdd
port 46 nsew
rlabel metal3 s 5668 11099 5766 11197 4 vdd
port 46 nsew
rlabel metal3 s 19227 11131 19325 11229 4 vdd
port 46 nsew
rlabel metal3 s 12939 4903 13037 5001 4 vdd
port 46 nsew
rlabel metal3 s 18427 14450 18525 14548 4 vdd
port 46 nsew
rlabel metal3 s 21565 9131 21663 9229 4 vdd
port 46 nsew
rlabel metal3 s 2555 9131 2653 9229 4 vdd
port 46 nsew
rlabel metal3 s 19227 11921 19325 12019 4 vdd
port 46 nsew
rlabel metal3 s 12253 6787 12351 6885 4 vdd
port 46 nsew
rlabel metal3 s 11748 7378 11846 7476 4 vdd
port 46 nsew
rlabel metal3 s 22888 8334 22986 8432 4 vdd
port 46 nsew
rlabel metal3 s 12441 4065 12539 4163 4 vdd
port 46 nsew
rlabel metal3 s 18452 8729 18550 8827 4 vdd
port 46 nsew
rlabel metal3 s 9757 15411 9855 15509 4 vdd
port 46 nsew
rlabel metal3 s 5668 8334 5766 8432 4 vdd
port 46 nsew
rlabel metal3 s 13620 7378 13718 7476 4 vdd
port 46 nsew
rlabel metal3 s 12253 15411 12351 15509 4 vdd
port 46 nsew
rlabel metal3 s 5668 10704 5766 10802 4 vdd
port 46 nsew
rlabel metal3 s 9933 4903 10031 5001 4 vdd
port 46 nsew
rlabel metal3 s 13501 15411 13599 15509 4 vdd
port 46 nsew
rlabel metal3 s 4893 13871 4991 13969 4 vdd
port 46 nsew
rlabel metal3 s 11124 14820 11222 14918 4 vdd
port 46 nsew
rlabel metal3 s 7564 7742 7662 7840 4 vdd
port 46 nsew
rlabel metal3 s 1232 10704 1330 10802 4 vdd
port 46 nsew
rlabel metal3 s 13677 17295 13775 17393 4 vdd
port 46 nsew
rlabel metal3 s 14175 18133 14273 18231 4 vdd
port 46 nsew
rlabel metal3 s 5668 12284 5766 12382 4 vdd
port 46 nsew
rlabel metal3 s 19227 12291 19325 12389 4 vdd
port 46 nsew
rlabel metal3 s 19227 13871 19325 13969 4 vdd
port 46 nsew
rlabel metal3 s 12927 4065 13025 4163 4 vdd
port 46 nsew
rlabel metal3 s 5668 12679 5766 12777 4 vdd
port 46 nsew
rlabel metal3 s 20790 10704 20888 10802 4 vdd
port 46 nsew
rlabel metal3 s 19227 9921 19325 10019 4 vdd
port 46 nsew
rlabel metal3 s 6525 7754 6623 7852 4 vdd
port 46 nsew
rlabel metal3 s 11193 18133 11291 18231 4 vdd
port 46 nsew
rlabel metal3 s 13584 1563 13682 1661 4 vdd
port 46 nsew
rlabel metal3 s 10431 3743 10529 3841 4 gnd
port 47 nsew
rlabel metal3 s 12511 16521 12609 16619 4 gnd
port 47 nsew
rlabel metal3 s 18848 9519 18946 9617 4 gnd
port 47 nsew
rlabel metal3 s 19652 13081 19750 13179 4 gnd
port 47 nsew
rlabel metal3 s 18020 11084 18118 11182 4 gnd
port 47 nsew
rlabel metal3 s 15564 9282 15662 9380 4 gnd
port 47 nsew
rlabel metal3 s 18848 12679 18946 12777 4 gnd
port 47 nsew
rlabel metal3 s 8556 10862 8654 10960 4 gnd
port 47 nsew
rlabel metal3 s 15564 8492 15662 8590 4 gnd
port 47 nsew
rlabel metal3 s 836 10704 934 10802 4 gnd
port 47 nsew
rlabel metal3 s 10015 16521 10113 16619 4 gnd
port 47 nsew
rlabel metal3 s 14175 3743 14273 3841 4 gnd
port 47 nsew
rlabel metal3 s 21990 10711 22088 10809 4 gnd
port 47 nsew
rlabel metal3 s 19652 11919 19750 12017 4 gnd
port 47 nsew
rlabel metal3 s 8556 8492 8654 8590 4 gnd
port 47 nsew
rlabel metal3 s 2934 10704 3032 10802 4 gnd
port 47 nsew
rlabel metal3 s 5272 8334 5370 8432 4 gnd
port 47 nsew
rlabel metal3 s 15564 8729 15662 8827 4 gnd
port 47 nsew
rlabel metal3 s 5272 9914 5370 10012 4 gnd
port 47 nsew
rlabel metal3 s 21990 9131 22088 9229 4 gnd
port 47 nsew
rlabel metal3 s 10361 5677 10459 5775 4 gnd
port 47 nsew
rlabel metal3 s 14165 2950 14263 3048 4 gnd
port 47 nsew
rlabel metal3 s 5272 13469 5370 13567 4 gnd
port 47 nsew
rlabel metal3 s 18848 11889 18946 11987 4 gnd
port 47 nsew
rlabel metal3 s 15564 9519 15662 9617 4 gnd
port 47 nsew
rlabel metal3 s 15564 8176 15662 8274 4 gnd
port 47 nsew
rlabel metal3 s 8556 8966 8654 9064 4 gnd
port 47 nsew
rlabel metal3 s 15564 8966 15662 9064 4 gnd
port 47 nsew
rlabel metal3 s 11679 3743 11777 3841 4 gnd
port 47 nsew
rlabel metal3 s 4468 13499 4566 13597 4 gnd
port 47 nsew
rlabel metal3 s 2934 8334 3032 8432 4 gnd
port 47 nsew
rlabel metal3 s 5272 11494 5370 11592 4 gnd
port 47 nsew
rlabel metal3 s 13689 18455 13787 18553 4 gnd
port 47 nsew
rlabel metal3 s 19652 13871 19750 13969 4 gnd
port 47 nsew
rlabel metal3 s 15564 12916 15662 13014 4 gnd
port 47 nsew
rlabel metal3 s 2130 11501 2228 11599 4 gnd
port 47 nsew
rlabel metal3 s 5272 12679 5370 12777 4 gnd
port 47 nsew
rlabel metal3 s 13570 1979 13668 2077 4 gnd
port 47 nsew
rlabel metal3 s 12807 2181 12905 2279 4 gnd
port 47 nsew
rlabel metal3 s 4468 10339 4566 10437 4 gnd
port 47 nsew
rlabel metal3 s 14105 5677 14203 5775 4 gnd
port 47 nsew
rlabel metal3 s 4468 9921 4566 10019 4 gnd
port 47 nsew
rlabel metal3 s 8190 7812 8288 7910 4 gnd
port 47 nsew
rlabel metal3 s 11609 5677 11707 5775 4 gnd
port 47 nsew
rlabel metal3 s 12511 5677 12609 5775 4 gnd
port 47 nsew
rlabel metal3 s 18848 9124 18946 9222 4 gnd
port 47 nsew
rlabel metal3 s 9826 1979 9924 2077 4 gnd
port 47 nsew
rlabel metal3 s 15564 10309 15662 10407 4 gnd
port 47 nsew
rlabel metal3 s 5272 9124 5370 9222 4 gnd
port 47 nsew
rlabel metal3 s 4468 13081 4566 13179 4 gnd
port 47 nsew
rlabel metal3 s 8190 0 8288 98 4 gnd
port 47 nsew
rlabel metal3 s 18848 11494 18946 11592 4 gnd
port 47 nsew
rlabel metal3 s 21990 11501 22088 11599 4 gnd
port 47 nsew
rlabel metal3 s 5272 8729 5370 8827 4 gnd
port 47 nsew
rlabel metal3 s 6100 11084 6198 11182 4 gnd
port 47 nsew
rlabel metal3 s 5272 11099 5370 11197 4 gnd
port 47 nsew
rlabel metal3 s 19652 9131 19750 9229 4 gnd
port 47 nsew
rlabel metal3 s 2130 8341 2228 8439 4 gnd
port 47 nsew
rlabel metal3 s 4468 8341 4566 8439 4 gnd
port 47 nsew
rlabel metal3 s 10431 18455 10529 18553 4 gnd
port 47 nsew
rlabel metal3 s 15564 11336 15662 11434 4 gnd
port 47 nsew
rlabel metal3 s 11189 2181 11287 2279 4 gnd
port 47 nsew
rlabel metal3 s 8556 14259 8654 14357 4 gnd
port 47 nsew
rlabel metal3 s 11074 1979 11172 2077 4 gnd
port 47 nsew
rlabel metal3 s 11079 2950 11177 3048 4 gnd
port 47 nsew
rlabel metal3 s 5272 10704 5370 10802 4 gnd
port 47 nsew
rlabel metal3 s 8556 9519 8654 9617 4 gnd
port 47 nsew
rlabel metal3 s 8556 8176 8654 8274 4 gnd
port 47 nsew
rlabel metal3 s 15564 12126 15662 12224 4 gnd
port 47 nsew
rlabel metal3 s 13685 2181 13783 2279 4 gnd
port 47 nsew
rlabel metal3 s 11609 16521 11707 16619 4 gnd
port 47 nsew
rlabel metal3 s 836 8334 934 8432 4 gnd
port 47 nsew
rlabel metal3 s 15564 10862 15662 10960 4 gnd
port 47 nsew
rlabel metal3 s 11669 2950 11767 3048 4 gnd
port 47 nsew
rlabel metal3 s 12857 5677 12955 5775 4 gnd
port 47 nsew
rlabel metal3 s 10426 1979 10524 2077 4 gnd
port 47 nsew
rlabel metal3 s 5272 13864 5370 13962 4 gnd
port 47 nsew
rlabel metal3 s 12441 18455 12539 18553 4 gnd
port 47 nsew
rlabel metal3 s 18848 13864 18946 13962 4 gnd
port 47 nsew
rlabel metal3 s 8556 14022 8654 14120 4 gnd
port 47 nsew
rlabel metal3 s 4468 12291 4566 12389 4 gnd
port 47 nsew
rlabel metal3 s 21990 8341 22088 8439 4 gnd
port 47 nsew
rlabel metal3 s 8556 7939 8654 8037 4 gnd
port 47 nsew
rlabel metal3 s 4468 12709 4566 12807 4 gnd
port 47 nsew
rlabel metal3 s 4468 11501 4566 11599 4 gnd
port 47 nsew
rlabel metal3 s 15564 14259 15662 14357 4 gnd
port 47 nsew
rlabel metal3 s 19652 9921 19750 10019 4 gnd
port 47 nsew
rlabel metal3 s 15930 7812 16028 7910 4 gnd
port 47 nsew
rlabel metal3 s 6942 11099 7040 11197 4 gnd
port 47 nsew
rlabel metal3 s 19652 8759 19750 8857 4 gnd
port 47 nsew
rlabel metal3 s 15564 11889 15662 11987 4 gnd
port 47 nsew
rlabel metal3 s 11674 1979 11772 2077 4 gnd
port 47 nsew
rlabel metal3 s 14175 18455 14273 18553 4 gnd
port 47 nsew
rlabel metal3 s 12917 2950 13015 3048 4 gnd
port 47 nsew
rlabel metal3 s 19652 9549 19750 9647 4 gnd
port 47 nsew
rlabel metal3 s 11193 18455 11291 18553 4 gnd
port 47 nsew
rlabel metal3 s 8556 11652 8654 11750 4 gnd
port 47 nsew
rlabel metal3 s 2934 11494 3032 11592 4 gnd
port 47 nsew
rlabel metal3 s 4468 11129 4566 11227 4 gnd
port 47 nsew
rlabel metal3 s 21186 8334 21284 8432 4 gnd
port 47 nsew
rlabel metal3 s 21186 9124 21284 9222 4 gnd
port 47 nsew
rlabel metal3 s 8190 14606 8288 14704 4 gnd
port 47 nsew
rlabel metal3 s 8556 9756 8654 9854 4 gnd
port 47 nsew
rlabel metal3 s 4468 9131 4566 9229 4 gnd
port 47 nsew
rlabel metal3 s 12441 3743 12539 3841 4 gnd
port 47 nsew
rlabel metal3 s 14055 2181 14153 2279 4 gnd
port 47 nsew
rlabel metal3 s 12857 16521 12955 16619 4 gnd
port 47 nsew
rlabel metal3 s 4468 10711 4566 10809 4 gnd
port 47 nsew
rlabel metal3 s 8556 12916 8654 13014 4 gnd
port 47 nsew
rlabel metal3 s 4468 13871 4566 13969 4 gnd
port 47 nsew
rlabel metal3 s 9945 18455 10043 18553 4 gnd
port 47 nsew
rlabel metal3 s 8556 13469 8654 13567 4 gnd
port 47 nsew
rlabel metal3 s 10015 5677 10113 5775 4 gnd
port 47 nsew
rlabel metal3 s 13759 16521 13857 16619 4 gnd
port 47 nsew
rlabel metal3 s 14170 1979 14268 2077 4 gnd
port 47 nsew
rlabel metal3 s 11263 16521 11361 16619 4 gnd
port 47 nsew
rlabel metal3 s 15564 13706 15662 13804 4 gnd
port 47 nsew
rlabel metal3 s 17178 11099 17276 11197 4 gnd
port 47 nsew
rlabel metal3 s 8556 12442 8654 12540 4 gnd
port 47 nsew
rlabel metal3 s 10361 16521 10459 16619 4 gnd
port 47 nsew
rlabel metal3 s 2934 9124 3032 9222 4 gnd
port 47 nsew
rlabel metal3 s 18848 10309 18946 10407 4 gnd
port 47 nsew
rlabel metal3 s 15564 10546 15662 10644 4 gnd
port 47 nsew
rlabel metal3 s 10421 2950 10519 3048 4 gnd
port 47 nsew
rlabel metal3 s 15564 13469 15662 13567 4 gnd
port 47 nsew
rlabel metal3 s 15930 14606 16028 14704 4 gnd
port 47 nsew
rlabel metal3 s 5272 12284 5370 12382 4 gnd
port 47 nsew
rlabel metal3 s 5272 11889 5370 11987 4 gnd
port 47 nsew
rlabel metal3 s 19652 13499 19750 13597 4 gnd
port 47 nsew
rlabel metal3 s 19652 12709 19750 12807 4 gnd
port 47 nsew
rlabel metal3 s 9945 3743 10043 3841 4 gnd
port 47 nsew
rlabel metal3 s 23284 10704 23382 10802 4 gnd
port 47 nsew
rlabel metal3 s 15564 12442 15662 12540 4 gnd
port 47 nsew
rlabel metal3 s 15564 9756 15662 9854 4 gnd
port 47 nsew
rlabel metal3 s 18848 8334 18946 8432 4 gnd
port 47 nsew
rlabel metal3 s 8556 10546 8654 10644 4 gnd
port 47 nsew
rlabel metal3 s 14556 0 14654 98 4 gnd
port 47 nsew
rlabel metal3 s 13759 5677 13857 5775 4 gnd
port 47 nsew
rlabel metal3 s 9831 2950 9929 3048 4 gnd
port 47 nsew
rlabel metal3 s 2130 9131 2228 9229 4 gnd
port 47 nsew
rlabel metal3 s 4468 8759 4566 8857 4 gnd
port 47 nsew
rlabel metal3 s 18848 12284 18946 12382 4 gnd
port 47 nsew
rlabel metal3 s 12322 1979 12420 2077 4 gnd
port 47 nsew
rlabel metal3 s 19652 12291 19750 12389 4 gnd
port 47 nsew
rlabel metal3 s 18848 9914 18946 10012 4 gnd
port 47 nsew
rlabel metal3 s 8556 13232 8654 13330 4 gnd
port 47 nsew
rlabel metal3 s 21186 11494 21284 11592 4 gnd
port 47 nsew
rlabel metal3 s 14105 16521 14203 16619 4 gnd
port 47 nsew
rlabel metal3 s 12437 2181 12535 2279 4 gnd
port 47 nsew
rlabel metal3 s 8556 8729 8654 8827 4 gnd
port 47 nsew
rlabel metal3 s 4468 11919 4566 12017 4 gnd
port 47 nsew
rlabel metal3 s 8556 11889 8654 11987 4 gnd
port 47 nsew
rlabel metal3 s 15564 14022 15662 14120 4 gnd
port 47 nsew
rlabel metal3 s 18848 10704 18946 10802 4 gnd
port 47 nsew
rlabel metal3 s 18848 8729 18946 8827 4 gnd
port 47 nsew
rlabel metal3 s 8556 13706 8654 13804 4 gnd
port 47 nsew
rlabel metal3 s 12927 3743 13025 3841 4 gnd
port 47 nsew
rlabel metal3 s 18848 13469 18946 13567 4 gnd
port 47 nsew
rlabel metal3 s 12922 1979 13020 2077 4 gnd
port 47 nsew
rlabel metal3 s 15564 12679 15662 12777 4 gnd
port 47 nsew
rlabel metal3 s 5272 9519 5370 9617 4 gnd
port 47 nsew
rlabel metal3 s 19652 11129 19750 11227 4 gnd
port 47 nsew
rlabel metal3 s 4468 9549 4566 9647 4 gnd
port 47 nsew
rlabel metal3 s 8556 12126 8654 12224 4 gnd
port 47 nsew
rlabel metal3 s 12927 18455 13025 18553 4 gnd
port 47 nsew
rlabel metal3 s 11559 2181 11657 2279 4 gnd
port 47 nsew
rlabel metal3 s 8556 10309 8654 10407 4 gnd
port 47 nsew
rlabel metal3 s 9941 2181 10039 2279 4 gnd
port 47 nsew
rlabel metal3 s 19652 8341 19750 8439 4 gnd
port 47 nsew
rlabel metal3 s 8556 12679 8654 12777 4 gnd
port 47 nsew
rlabel metal3 s 15564 11652 15662 11750 4 gnd
port 47 nsew
rlabel metal3 s 5272 13074 5370 13172 4 gnd
port 47 nsew
rlabel metal3 s 19652 10339 19750 10437 4 gnd
port 47 nsew
rlabel metal3 s 8556 9282 8654 9380 4 gnd
port 47 nsew
rlabel metal3 s 13689 3743 13787 3841 4 gnd
port 47 nsew
rlabel metal3 s 8556 11336 8654 11434 4 gnd
port 47 nsew
rlabel metal3 s 5272 10309 5370 10407 4 gnd
port 47 nsew
rlabel metal3 s 19652 10711 19750 10809 4 gnd
port 47 nsew
rlabel metal3 s 15564 10072 15662 10170 4 gnd
port 47 nsew
rlabel metal3 s 8556 11099 8654 11197 4 gnd
port 47 nsew
rlabel metal3 s 21186 10704 21284 10802 4 gnd
port 47 nsew
rlabel metal3 s 18848 11099 18946 11197 4 gnd
port 47 nsew
rlabel metal3 s 19652 11501 19750 11599 4 gnd
port 47 nsew
rlabel metal3 s 11263 5677 11361 5775 4 gnd
port 47 nsew
rlabel metal3 s 23284 8334 23382 8432 4 gnd
port 47 nsew
rlabel metal3 s 15564 7939 15662 8037 4 gnd
port 47 nsew
rlabel metal3 s 18848 13074 18946 13172 4 gnd
port 47 nsew
rlabel metal3 s 11679 18455 11777 18553 4 gnd
port 47 nsew
rlabel metal3 s 15564 11099 15662 11197 4 gnd
port 47 nsew
rlabel metal3 s 10311 2181 10409 2279 4 gnd
port 47 nsew
rlabel metal3 s 2130 10711 2228 10809 4 gnd
port 47 nsew
rlabel metal3 s 11193 3743 11291 3841 4 gnd
port 47 nsew
rlabel metal3 s 12327 2950 12425 3048 4 gnd
port 47 nsew
rlabel metal3 s 8556 10072 8654 10170 4 gnd
port 47 nsew
rlabel metal3 s 13575 2950 13673 3048 4 gnd
port 47 nsew
rlabel metal3 s 15564 13232 15662 13330 4 gnd
port 47 nsew
<< properties >>
string FIXED_BBOX 0 0 24302 18647
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 462292
string GDS_START 362780
<< end >>
