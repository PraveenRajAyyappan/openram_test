magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1335 -1309 7878 19691
<< locali >>
rect 6517 8501 6551 8517
rect 4178 8467 6517 8501
rect 6517 8451 6551 8467
rect 3290 7832 3324 7848
rect 3290 7782 3324 7798
rect 3883 7794 3917 7810
rect 3883 7744 3917 7760
rect 6517 7087 6551 7103
rect 4178 7053 6517 7087
rect 6517 7037 6551 7053
rect 3573 6790 3792 6824
rect 3758 6308 3792 6790
rect 4245 6343 4279 6359
rect 4245 6293 4279 6309
rect 3438 6191 3472 6207
rect 3438 6141 3472 6157
rect 3338 5943 3372 5959
rect 3338 5893 3372 5909
rect 6517 5673 6551 5689
rect 4504 5639 6517 5673
rect 6517 5623 6551 5639
rect 3305 5403 3339 5419
rect 3305 5353 3339 5369
rect 3438 5279 3472 5295
rect 3438 5229 3472 5245
rect 3571 5155 3605 5171
rect 3571 5105 3605 5121
rect 4101 4982 4135 4998
rect 4101 4932 4135 4948
rect 6517 4259 6551 4275
rect 4504 4225 6517 4259
rect 6517 4209 6551 4225
rect 4109 3536 4143 3552
rect 4109 3486 4143 3502
rect 3438 3363 3472 3379
rect 3438 3313 3472 3329
rect 3338 3115 3372 3131
rect 3338 3065 3372 3081
rect 6517 2845 6551 2861
rect 4620 2811 6517 2845
rect 6517 2795 6551 2811
rect 3555 2541 3740 2575
rect 3290 2176 3324 2192
rect 3555 2176 3589 2541
rect 3806 2327 3840 2343
rect 3806 2277 3840 2293
rect 3422 2142 3589 2176
rect 4477 2154 4511 2170
rect 3290 2126 3324 2142
rect 4477 2104 4511 2120
rect 6517 1431 6551 1447
rect 4988 1397 6517 1431
rect 6517 1381 6551 1397
rect 5699 724 5733 740
rect 3290 686 3324 702
rect 5699 674 5733 690
rect 3290 636 3324 652
rect 6517 17 6551 33
rect 6517 -33 6551 -17
<< viali >>
rect 6517 8467 6551 8501
rect 3290 7798 3324 7832
rect 3883 7760 3917 7794
rect 6517 7053 6551 7087
rect 4245 6309 4279 6343
rect 3438 6157 3472 6191
rect 3338 5909 3372 5943
rect 6517 5639 6551 5673
rect 3305 5369 3339 5403
rect 3438 5245 3472 5279
rect 3571 5121 3605 5155
rect 4101 4948 4135 4982
rect 6517 4225 6551 4259
rect 4109 3502 4143 3536
rect 3438 3329 3472 3363
rect 3338 3081 3372 3115
rect 6517 2811 6551 2845
rect 3806 2293 3840 2327
rect 3290 2142 3324 2176
rect 4477 2120 4511 2154
rect 6517 1397 6551 1431
rect 3290 652 3324 686
rect 5699 690 5733 724
rect 6517 -17 6551 17
<< metal1 >>
rect 6502 8458 6508 8510
rect 6560 8458 6566 8510
rect 2704 7789 2710 7841
rect 2762 7829 2768 7841
rect 3278 7832 3336 7838
rect 3278 7829 3290 7832
rect 2762 7801 3290 7829
rect 2762 7789 2768 7801
rect 3278 7798 3290 7801
rect 3324 7798 3336 7832
rect 3278 7792 3336 7798
rect 3868 7751 3874 7803
rect 3926 7751 3932 7803
rect 6502 7044 6508 7096
rect 6560 7044 6566 7096
rect 4230 6300 4236 6352
rect 4288 6300 4294 6352
rect 2620 6148 2626 6200
rect 2678 6188 2684 6200
rect 3426 6191 3484 6197
rect 3426 6188 3438 6191
rect 2678 6160 3438 6188
rect 2678 6148 2684 6160
rect 3426 6157 3438 6160
rect 3472 6157 3484 6191
rect 3426 6151 3484 6157
rect 2788 5900 2794 5952
rect 2846 5940 2852 5952
rect 3326 5943 3384 5949
rect 3326 5940 3338 5943
rect 2846 5912 3338 5940
rect 2846 5900 2852 5912
rect 3326 5909 3338 5912
rect 3372 5909 3384 5943
rect 3326 5903 3384 5909
rect 6502 5630 6508 5682
rect 6560 5630 6566 5682
rect 2620 5360 2626 5412
rect 2678 5400 2684 5412
rect 3293 5403 3351 5409
rect 3293 5400 3305 5403
rect 2678 5372 3305 5400
rect 2678 5360 2684 5372
rect 3293 5369 3305 5372
rect 3339 5369 3351 5403
rect 3293 5363 3351 5369
rect 2704 5236 2710 5288
rect 2762 5276 2768 5288
rect 3426 5279 3484 5285
rect 3426 5276 3438 5279
rect 2762 5248 3438 5276
rect 2762 5236 2768 5248
rect 3426 5245 3438 5248
rect 3472 5245 3484 5279
rect 3426 5239 3484 5245
rect 3040 5112 3046 5164
rect 3098 5152 3104 5164
rect 3559 5155 3617 5161
rect 3559 5152 3571 5155
rect 3098 5124 3571 5152
rect 3098 5112 3104 5124
rect 3559 5121 3571 5124
rect 3605 5121 3617 5155
rect 3559 5115 3617 5121
rect 4086 4939 4092 4991
rect 4144 4939 4150 4991
rect 1521 4296 1527 4348
rect 1579 4336 1585 4348
rect 2620 4336 2626 4348
rect 1579 4308 2626 4336
rect 1579 4296 1585 4308
rect 2620 4296 2626 4308
rect 2678 4296 2684 4348
rect 6502 4216 6508 4268
rect 6560 4216 6566 4268
rect 351 4136 357 4188
rect 409 4176 415 4188
rect 2872 4176 2878 4188
rect 409 4148 2878 4176
rect 409 4136 415 4148
rect 2872 4136 2878 4148
rect 2930 4136 2936 4188
rect 4094 3493 4100 3545
rect 4152 3493 4158 3545
rect 3040 3320 3046 3372
rect 3098 3360 3104 3372
rect 3426 3363 3484 3369
rect 3426 3360 3438 3363
rect 3098 3332 3438 3360
rect 3098 3320 3104 3332
rect 3426 3329 3438 3332
rect 3472 3329 3484 3363
rect 3426 3323 3484 3329
rect 2872 3072 2878 3124
rect 2930 3112 2936 3124
rect 3326 3115 3384 3121
rect 3326 3112 3338 3115
rect 2930 3084 3338 3112
rect 2930 3072 2936 3084
rect 3326 3081 3338 3084
rect 3372 3081 3384 3115
rect 3326 3075 3384 3081
rect 6502 2802 6508 2854
rect 6560 2802 6566 2854
rect 3791 2284 3797 2336
rect 3849 2284 3855 2336
rect 2872 2133 2878 2185
rect 2930 2173 2936 2185
rect 3278 2176 3336 2182
rect 3278 2173 3290 2176
rect 2930 2145 3290 2173
rect 2930 2133 2936 2145
rect 3278 2142 3290 2145
rect 3324 2142 3336 2176
rect 3278 2136 3336 2142
rect 4462 2111 4468 2163
rect 4520 2111 4526 2163
rect 6502 1388 6508 1440
rect 6560 1388 6566 1440
rect 3275 643 3281 695
rect 3333 643 3339 695
rect 5684 681 5690 733
rect 5742 681 5748 733
rect 6502 -26 6508 26
rect 6560 -26 6566 26
<< via1 >>
rect 6508 8501 6560 8510
rect 6508 8467 6517 8501
rect 6517 8467 6551 8501
rect 6551 8467 6560 8501
rect 6508 8458 6560 8467
rect 2710 7789 2762 7841
rect 3874 7794 3926 7803
rect 3874 7760 3883 7794
rect 3883 7760 3917 7794
rect 3917 7760 3926 7794
rect 3874 7751 3926 7760
rect 6508 7087 6560 7096
rect 6508 7053 6517 7087
rect 6517 7053 6551 7087
rect 6551 7053 6560 7087
rect 6508 7044 6560 7053
rect 4236 6343 4288 6352
rect 4236 6309 4245 6343
rect 4245 6309 4279 6343
rect 4279 6309 4288 6343
rect 4236 6300 4288 6309
rect 2626 6148 2678 6200
rect 2794 5900 2846 5952
rect 6508 5673 6560 5682
rect 6508 5639 6517 5673
rect 6517 5639 6551 5673
rect 6551 5639 6560 5673
rect 6508 5630 6560 5639
rect 2626 5360 2678 5412
rect 2710 5236 2762 5288
rect 3046 5112 3098 5164
rect 4092 4982 4144 4991
rect 4092 4948 4101 4982
rect 4101 4948 4135 4982
rect 4135 4948 4144 4982
rect 4092 4939 4144 4948
rect 1527 4296 1579 4348
rect 2626 4296 2678 4348
rect 6508 4259 6560 4268
rect 6508 4225 6517 4259
rect 6517 4225 6551 4259
rect 6551 4225 6560 4259
rect 6508 4216 6560 4225
rect 357 4136 409 4188
rect 2878 4136 2930 4188
rect 4100 3536 4152 3545
rect 4100 3502 4109 3536
rect 4109 3502 4143 3536
rect 4143 3502 4152 3536
rect 4100 3493 4152 3502
rect 3046 3320 3098 3372
rect 2878 3072 2930 3124
rect 6508 2845 6560 2854
rect 6508 2811 6517 2845
rect 6517 2811 6551 2845
rect 6551 2811 6560 2845
rect 6508 2802 6560 2811
rect 3797 2327 3849 2336
rect 3797 2293 3806 2327
rect 3806 2293 3840 2327
rect 3840 2293 3849 2327
rect 3797 2284 3849 2293
rect 2878 2133 2930 2185
rect 4468 2154 4520 2163
rect 4468 2120 4477 2154
rect 4477 2120 4511 2154
rect 4511 2120 4520 2154
rect 4468 2111 4520 2120
rect 6508 1431 6560 1440
rect 6508 1397 6517 1431
rect 6517 1397 6551 1431
rect 6551 1397 6560 1431
rect 6508 1388 6560 1397
rect 3281 686 3333 695
rect 3281 652 3290 686
rect 3290 652 3324 686
rect 3324 652 3333 686
rect 3281 643 3333 652
rect 5690 724 5742 733
rect 5690 690 5699 724
rect 5699 690 5733 724
rect 5733 690 5742 724
rect 5690 681 5742 690
rect 6508 17 6560 26
rect 6508 -17 6517 17
rect 6517 -17 6551 17
rect 6551 -17 6560 17
rect 6508 -26 6560 -17
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4354 1567 6401
rect 1527 4348 1579 4354
rect 1527 4290 1579 4296
rect 357 4188 409 4194
rect 357 4130 409 4136
rect 369 1414 397 4130
rect 1844 913 1900 922
rect 1844 848 1900 857
rect 137 538 203 590
rect 2350 531 2406 540
rect 2350 466 2406 475
rect 2554 0 2582 8524
rect 2638 6206 2666 8524
rect 2722 7847 2750 8524
rect 2710 7841 2762 7847
rect 2710 7783 2762 7789
rect 2626 6200 2678 6206
rect 2626 6142 2678 6148
rect 2638 5418 2666 6142
rect 2626 5412 2678 5418
rect 2626 5354 2678 5360
rect 2638 4354 2666 5354
rect 2722 5294 2750 7783
rect 2806 5958 2834 8524
rect 2794 5952 2846 5958
rect 2794 5894 2846 5900
rect 2710 5288 2762 5294
rect 2710 5230 2762 5236
rect 2626 4348 2678 4354
rect 2626 4290 2678 4296
rect 2638 0 2666 4290
rect 2722 1608 2750 5230
rect 2806 3556 2834 5894
rect 2890 4194 2918 8524
rect 2878 4188 2930 4194
rect 2878 4130 2930 4136
rect 2792 3547 2848 3556
rect 2792 3482 2848 3491
rect 2708 1599 2764 1608
rect 2708 1534 2764 1543
rect 2722 0 2750 1534
rect 2806 0 2834 3482
rect 2890 3130 2918 4130
rect 2878 3124 2930 3130
rect 2878 3066 2930 3072
rect 2890 2191 2918 3066
rect 2878 2185 2930 2191
rect 2878 2127 2930 2133
rect 2890 178 2918 2127
rect 2974 540 3002 8524
rect 3058 5170 3086 8524
rect 6506 8512 6562 8521
rect 6506 8447 6562 8456
rect 3874 7803 3926 7809
rect 3926 7763 6618 7791
rect 3874 7745 3926 7751
rect 6506 7098 6562 7107
rect 6506 7033 6562 7042
rect 4236 6352 4288 6358
rect 4288 6312 6618 6340
rect 4236 6294 4288 6300
rect 6506 5684 6562 5693
rect 6506 5619 6562 5628
rect 3046 5164 3098 5170
rect 3046 5106 3098 5112
rect 3058 3378 3086 5106
rect 4092 4991 4144 4997
rect 4144 4951 6618 4979
rect 4092 4933 4144 4939
rect 6506 4270 6562 4279
rect 6506 4205 6562 4214
rect 4098 3547 4154 3556
rect 4098 3482 4154 3491
rect 3046 3372 3098 3378
rect 3046 3314 3098 3320
rect 3058 2347 3086 3314
rect 6506 2856 6562 2865
rect 6506 2791 6562 2800
rect 3044 2338 3100 2347
rect 3044 2273 3100 2282
rect 3795 2338 3851 2347
rect 3795 2273 3851 2282
rect 3058 922 3086 2273
rect 4468 2163 4520 2169
rect 4468 2105 4520 2111
rect 4480 1608 4508 2105
rect 4466 1599 4522 1608
rect 4466 1534 4522 1543
rect 6506 1442 6562 1451
rect 6506 1377 6562 1386
rect 3044 913 3100 922
rect 3044 848 3100 857
rect 2960 531 3016 540
rect 2960 466 3016 475
rect 2876 169 2932 178
rect 2876 104 2932 113
rect 2890 0 2918 104
rect 2974 0 3002 466
rect 3058 0 3086 848
rect 5690 733 5742 739
rect 3281 695 3333 701
rect 5742 693 6618 721
rect 5690 675 5742 681
rect 3281 637 3333 643
rect 5702 178 5730 675
rect 5688 169 5744 178
rect 5688 104 5744 113
rect 6506 28 6562 37
rect 6506 -37 6562 -28
<< via2 >>
rect 1844 857 1900 913
rect 2350 475 2406 531
rect 2792 3491 2848 3547
rect 2708 1543 2764 1599
rect 6506 8510 6562 8512
rect 6506 8458 6508 8510
rect 6508 8458 6560 8510
rect 6560 8458 6562 8510
rect 6506 8456 6562 8458
rect 6506 7096 6562 7098
rect 6506 7044 6508 7096
rect 6508 7044 6560 7096
rect 6560 7044 6562 7096
rect 6506 7042 6562 7044
rect 6506 5682 6562 5684
rect 6506 5630 6508 5682
rect 6508 5630 6560 5682
rect 6560 5630 6562 5682
rect 6506 5628 6562 5630
rect 6506 4268 6562 4270
rect 6506 4216 6508 4268
rect 6508 4216 6560 4268
rect 6560 4216 6562 4268
rect 6506 4214 6562 4216
rect 4098 3545 4154 3547
rect 4098 3493 4100 3545
rect 4100 3493 4152 3545
rect 4152 3493 4154 3545
rect 4098 3491 4154 3493
rect 6506 2854 6562 2856
rect 6506 2802 6508 2854
rect 6508 2802 6560 2854
rect 6560 2802 6562 2854
rect 6506 2800 6562 2802
rect 3044 2282 3100 2338
rect 3795 2336 3851 2338
rect 3795 2284 3797 2336
rect 3797 2284 3849 2336
rect 3849 2284 3851 2336
rect 3795 2282 3851 2284
rect 4466 1543 4522 1599
rect 6506 1440 6562 1442
rect 6506 1388 6508 1440
rect 6508 1388 6560 1440
rect 6560 1388 6562 1440
rect 6506 1386 6562 1388
rect 3044 857 3100 913
rect 2960 475 3016 531
rect 2876 113 2932 169
rect 5688 113 5744 169
rect 6506 26 6562 28
rect 6506 -26 6508 26
rect 6508 -26 6560 26
rect 6560 -26 6562 26
rect 6506 -28 6562 -26
<< metal3 >>
rect 607 18333 705 18431
rect 1343 18333 1441 18431
rect 607 16919 705 17017
rect 1343 16919 1441 17017
rect 607 15505 705 15603
rect 1343 15505 1441 15603
rect 607 14091 705 14189
rect 1343 14091 1441 14189
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 6485 8512 6583 8533
rect 6485 8456 6506 8512
rect 6562 8456 6583 8512
rect 6485 8435 6583 8456
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 6485 7098 6583 7119
rect 6485 7042 6506 7098
rect 6562 7042 6583 7098
rect 6485 7021 6583 7042
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 6485 5684 6583 5705
rect 6485 5628 6506 5684
rect 6562 5628 6583 5684
rect 6485 5607 6583 5628
rect 6485 4270 6583 4291
rect 6485 4214 6506 4270
rect 6562 4214 6583 4270
rect 6485 4193 6583 4214
rect 2787 3549 2853 3552
rect 4093 3549 4159 3552
rect 2787 3547 4159 3549
rect 2787 3491 2792 3547
rect 2848 3491 4098 3547
rect 4154 3491 4159 3547
rect 2787 3489 4159 3491
rect 2787 3486 2853 3489
rect 4093 3486 4159 3489
rect 6485 2856 6583 2877
rect 6485 2800 6506 2856
rect 6562 2800 6583 2856
rect 6485 2779 6583 2800
rect 3039 2340 3105 2343
rect 3790 2340 3856 2343
rect 3039 2338 3856 2340
rect 3039 2282 3044 2338
rect 3100 2282 3795 2338
rect 3851 2282 3856 2338
rect 3039 2280 3856 2282
rect 3039 2277 3105 2280
rect 3790 2277 3856 2280
rect 2703 1601 2769 1604
rect 4461 1601 4527 1604
rect 2703 1599 4527 1601
rect 2703 1543 2708 1599
rect 2764 1543 4466 1599
rect 4522 1543 4527 1599
rect 2703 1541 4527 1543
rect 2703 1538 2769 1541
rect 4461 1538 4527 1541
rect -49 1365 49 1463
rect 6485 1442 6583 1463
rect 6485 1386 6506 1442
rect 6562 1386 6583 1442
rect 6485 1365 6583 1386
rect 1839 915 1905 918
rect 3039 915 3105 918
rect 1839 913 3105 915
rect 1839 857 1844 913
rect 1900 857 3044 913
rect 3100 857 3105 913
rect 1839 855 3105 857
rect 1839 852 1905 855
rect 3039 852 3105 855
rect 2345 533 2411 536
rect 2955 533 3021 536
rect 2345 531 3021 533
rect 2345 475 2350 531
rect 2406 475 2960 531
rect 3016 475 3021 531
rect 2345 473 3021 475
rect 2345 470 2411 473
rect 2955 470 3021 473
rect 2871 171 2937 174
rect 5683 171 5749 174
rect 2871 169 5749 171
rect 2871 113 2876 169
rect 2932 113 5688 169
rect 5744 113 5749 169
rect 2871 111 5749 113
rect 2871 108 2937 111
rect 5683 108 5749 111
rect -49 -49 49 49
rect 6485 28 6583 49
rect 6485 -28 6506 28
rect 6562 -28 6583 28
rect 6485 -49 6583 -28
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 6501 0 1 8447
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 6502 0 1 8452
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 6505 0 1 8451
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 6501 0 1 7033
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 6502 0 1 7038
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 6505 0 1 7037
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 6501 0 1 5619
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 6502 0 1 5624
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 6505 0 1 5623
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 6501 0 1 7033
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 6502 0 1 7038
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 6505 0 1 7037
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 6501 0 1 5619
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 6502 0 1 5624
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 6505 0 1 5623
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 6501 0 1 4205
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 6502 0 1 4210
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 6505 0 1 4209
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 6501 0 1 2791
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 6502 0 1 2796
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 6505 0 1 2795
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 6501 0 1 4205
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 6502 0 1 4210
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 6505 0 1 4209
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 6501 0 1 2791
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 6502 0 1 2796
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 6505 0 1 2795
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 6501 0 1 1377
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 6502 0 1 1382
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 6505 0 1 1381
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 6501 0 1 -37
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 6502 0 1 -32
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 6505 0 1 -33
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 6501 0 1 1377
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 6502 0 1 1382
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 6505 0 1 1381
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 4094 0 1 3487
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1634918361
transform 1 0 4097 0 1 3486
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 4093 0 1 3482
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 4094 0 1 3487
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1634918361
transform 1 0 4097 0 1 3486
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1634918361
transform 1 0 2787 0 1 3482
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1634918361
transform 1 0 3426 0 1 3313
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 3040 0 1 3314
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1634918361
transform 1 0 3326 0 1 3065
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 2872 0 1 3066
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1634918361
transform 1 0 4462 0 1 2105
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1634918361
transform 1 0 4465 0 1 2104
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1634918361
transform 1 0 2703 0 1 1534
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1634918361
transform 1 0 4461 0 1 1534
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 3790 0 1 2273
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1634918361
transform 1 0 3791 0 1 2278
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1634918361
transform 1 0 3794 0 1 2277
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 3790 0 1 2273
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1634918361
transform 1 0 3791 0 1 2278
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1634918361
transform 1 0 3794 0 1 2277
box 0 0 1 1
use contact_29  contact_29_3
timestamp 1634918361
transform 1 0 3039 0 1 2273
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1634918361
transform 1 0 3278 0 1 2126
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1634918361
transform 1 0 2872 0 1 2127
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1634918361
transform 1 0 5684 0 1 675
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1634918361
transform 1 0 5687 0 1 674
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1634918361
transform 1 0 5684 0 1 675
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1634918361
transform 1 0 5687 0 1 674
box 0 0 1 1
use contact_29  contact_29_4
timestamp 1634918361
transform 1 0 2871 0 1 104
box 0 0 1 1
use contact_29  contact_29_5
timestamp 1634918361
transform 1 0 5683 0 1 104
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1634918361
transform 1 0 3275 0 1 637
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1634918361
transform 1 0 3278 0 1 636
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1634918361
transform 1 0 4230 0 1 6294
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1634918361
transform 1 0 4233 0 1 6293
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1634918361
transform 1 0 3426 0 1 6141
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1634918361
transform 1 0 2620 0 1 6142
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1634918361
transform 1 0 3326 0 1 5893
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1634918361
transform 1 0 2788 0 1 5894
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1634918361
transform 1 0 2620 0 1 4290
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1634918361
transform 1 0 1521 0 1 4290
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1634918361
transform 1 0 4086 0 1 4933
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1634918361
transform 1 0 4089 0 1 4932
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1634918361
transform 1 0 3559 0 1 5105
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1634918361
transform 1 0 3040 0 1 5106
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1634918361
transform 1 0 3426 0 1 5229
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1634918361
transform 1 0 2704 0 1 5230
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1634918361
transform 1 0 3293 0 1 5353
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1634918361
transform 1 0 2620 0 1 5354
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1634918361
transform 1 0 3868 0 1 7745
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1634918361
transform 1 0 3871 0 1 7744
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1634918361
transform 1 0 3278 0 1 7782
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1634918361
transform 1 0 2704 0 1 7783
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1634918361
transform 1 0 2872 0 1 4130
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1634918361
transform 1 0 351 0 1 4130
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 2345 0 1 466
box 0 0 1 1
use contact_29  contact_29_6
timestamp 1634918361
transform 1 0 2955 0 1 466
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 1839 0 1 848
box 0 0 1 1
use contact_29  contact_29_7
timestamp 1634918361
transform 1 0 3039 0 1 848
box 0 0 1 1
use pdriver_5  pdriver_5_0
timestamp 1634918361
transform 1 0 3694 0 1 5656
box -36 -17 880 1471
use pnand2_1  pnand2_1_0
timestamp 1634918361
transform 1 0 3226 0 1 5656
box -36 -17 504 1471
use delay_chain  delay_chain_0
timestamp 1634918361
transform 1 0 0 0 -1 18382
box -75 -49 1876 12783
use pand3_0  pand3_0_0
timestamp 1634918361
transform 1 0 3226 0 -1 5656
box -36 -17 1314 1471
use pdriver_2  pdriver_2_0
timestamp 1634918361
transform 1 0 3226 0 -1 8484
box -36 -17 988 1471
use pand2_0  pand2_0_0
timestamp 1634918361
transform 1 0 3226 0 1 2828
box -36 -17 1430 1471
use pand2_0  pand2_0_1
timestamp 1634918361
transform 1 0 3594 0 -1 2828
box -36 -17 1430 1471
use pinv_10  pinv_10_0
timestamp 1634918361
transform 1 0 3226 0 -1 2828
box -36 -17 404 1471
use pdriver_6  pdriver_6_0
timestamp 1634918361
transform 1 0 3226 0 1 0
box -36 -17 3344 1471
use dff_buf_array_0  dff_buf_array_0_0
timestamp 1634918361
transform 1 0 0 0 1 0
box -49 -49 2590 1471
<< labels >>
rlabel metal2 s 137 538 203 590 4 csb
port 1 nsew
rlabel metal2 s 3900 7763 6618 7791 4 wl_en
port 2 nsew
rlabel metal2 s 4118 4951 6618 4979 4 s_en
port 3 nsew
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
port 4 nsew
rlabel metal2 s 4262 6312 6618 6340 4 p_en_bar
port 5 nsew
rlabel metal2 s 3293 655 3321 683 4 clk
port 6 nsew
rlabel metal2 s 5716 693 6618 721 4 clk_buf
port 7 nsew
rlabel metal3 s 1343 5607 1441 5705 4 vdd
port 8 nsew
rlabel metal3 s 1343 11263 1441 11361 4 vdd
port 8 nsew
rlabel metal3 s 6485 4193 6583 4291 4 vdd
port 8 nsew
rlabel metal3 s 1343 14091 1441 14189 4 vdd
port 8 nsew
rlabel metal3 s 6485 1365 6583 1463 4 vdd
port 8 nsew
rlabel metal3 s 607 14091 705 14189 4 vdd
port 8 nsew
rlabel metal3 s 607 11263 705 11361 4 vdd
port 8 nsew
rlabel metal3 s 607 8435 705 8533 4 vdd
port 8 nsew
rlabel metal3 s 1343 16919 1441 17017 4 vdd
port 8 nsew
rlabel metal3 s 607 5607 705 5705 4 vdd
port 8 nsew
rlabel metal3 s 607 16919 705 17017 4 vdd
port 8 nsew
rlabel metal3 s -49 1365 49 1463 4 vdd
port 8 nsew
rlabel metal3 s 6485 7021 6583 7119 4 vdd
port 8 nsew
rlabel metal3 s 1343 8435 1441 8533 4 vdd
port 8 nsew
rlabel metal3 s 6485 5607 6583 5705 4 gnd
port 9 nsew
rlabel metal3 s 607 15505 705 15603 4 gnd
port 9 nsew
rlabel metal3 s 1343 15505 1441 15603 4 gnd
port 9 nsew
rlabel metal3 s 607 18333 705 18431 4 gnd
port 9 nsew
rlabel metal3 s 607 7021 705 7119 4 gnd
port 9 nsew
rlabel metal3 s 1343 18333 1441 18431 4 gnd
port 9 nsew
rlabel metal3 s 1343 9849 1441 9947 4 gnd
port 9 nsew
rlabel metal3 s -49 -49 49 49 4 gnd
port 9 nsew
rlabel metal3 s 6485 2779 6583 2877 4 gnd
port 9 nsew
rlabel metal3 s 607 9849 705 9947 4 gnd
port 9 nsew
rlabel metal3 s 6485 -49 6583 49 4 gnd
port 9 nsew
rlabel metal3 s 607 12677 705 12775 4 gnd
port 9 nsew
rlabel metal3 s 6485 8435 6583 8533 4 gnd
port 9 nsew
rlabel metal3 s 1343 7021 1441 7119 4 gnd
port 9 nsew
rlabel metal3 s 1343 12677 1441 12775 4 gnd
port 9 nsew
<< properties >>
string FIXED_BBOX 6501 -37 6567 0
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1194906
string GDS_START 1177916
<< end >>
