magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1260 -1260 8167 3516
<< metal1 >>
rect 1465 2168 1471 2220
rect 1523 2168 1529 2220
rect 1570 1130 1604 2256
rect 1646 1142 1674 2256
rect 1793 2016 1799 2068
rect 1851 2016 1857 2068
rect 2139 2016 2145 2068
rect 2197 2016 2203 2068
rect 1711 1242 1717 1294
rect 1769 1242 1775 1294
rect 2221 1242 2227 1294
rect 2279 1242 2285 1294
rect 2322 1142 2350 2256
rect 2392 1130 2426 2256
rect 2467 2168 2473 2220
rect 2525 2168 2531 2220
rect 2713 2168 2719 2220
rect 2771 2168 2777 2220
rect 2818 1130 2852 2256
rect 2894 1142 2922 2256
rect 3041 2016 3047 2068
rect 3099 2016 3105 2068
rect 3387 2016 3393 2068
rect 3445 2016 3451 2068
rect 2959 1242 2965 1294
rect 3017 1242 3023 1294
rect 3469 1242 3475 1294
rect 3527 1242 3533 1294
rect 3570 1142 3598 2256
rect 3640 1130 3674 2256
rect 3715 2168 3721 2220
rect 3773 2168 3779 2220
rect 3961 2168 3967 2220
rect 4019 2168 4025 2220
rect 4066 1130 4100 2256
rect 4142 1142 4170 2256
rect 4289 2016 4295 2068
rect 4347 2016 4353 2068
rect 4635 2016 4641 2068
rect 4693 2016 4699 2068
rect 4207 1242 4213 1294
rect 4265 1242 4271 1294
rect 4717 1242 4723 1294
rect 4775 1242 4781 1294
rect 4818 1142 4846 2256
rect 4888 1130 4922 2256
rect 4963 2168 4969 2220
rect 5021 2168 5027 2220
rect 5209 2168 5215 2220
rect 5267 2168 5273 2220
rect 5314 1130 5348 2256
rect 5390 1142 5418 2256
rect 5537 2016 5543 2068
rect 5595 2016 5601 2068
rect 5883 2016 5889 2068
rect 5941 2016 5947 2068
rect 5455 1242 5461 1294
rect 5513 1242 5519 1294
rect 5965 1242 5971 1294
rect 6023 1242 6029 1294
rect 6066 1142 6094 2256
rect 6136 1130 6170 2256
rect 6211 2168 6217 2220
rect 6269 2168 6275 2220
rect 1723 404 1729 456
rect 1781 404 1787 456
rect 2209 404 2215 456
rect 2267 404 2273 456
rect 2971 404 2977 456
rect 3029 404 3035 456
rect 3457 404 3463 456
rect 3515 404 3521 456
rect 4219 404 4225 456
rect 4277 404 4283 456
rect 4705 404 4711 456
rect 4763 404 4769 456
rect 5467 404 5473 456
rect 5525 404 5531 456
rect 5953 404 5959 456
rect 6011 404 6017 456
rect 1478 0 1524 254
rect 1723 82 1729 134
rect 1781 82 1787 134
rect 2209 82 2215 134
rect 2267 82 2273 134
rect 2472 0 2518 254
rect 2726 0 2772 254
rect 2971 82 2977 134
rect 3029 82 3035 134
rect 3457 82 3463 134
rect 3515 82 3521 134
rect 3720 0 3766 254
rect 3974 0 4020 254
rect 4219 82 4225 134
rect 4277 82 4283 134
rect 4705 82 4711 134
rect 4763 82 4769 134
rect 4968 0 5014 254
rect 5222 0 5268 254
rect 5467 82 5473 134
rect 5525 82 5531 134
rect 5953 82 5959 134
rect 6011 82 6017 134
rect 6216 0 6262 254
<< via1 >>
rect 1471 2168 1523 2220
rect 1799 2016 1851 2068
rect 2145 2016 2197 2068
rect 1717 1242 1769 1294
rect 2227 1242 2279 1294
rect 2473 2168 2525 2220
rect 2719 2168 2771 2220
rect 3047 2016 3099 2068
rect 3393 2016 3445 2068
rect 2965 1242 3017 1294
rect 3475 1242 3527 1294
rect 3721 2168 3773 2220
rect 3967 2168 4019 2220
rect 4295 2016 4347 2068
rect 4641 2016 4693 2068
rect 4213 1242 4265 1294
rect 4723 1242 4775 1294
rect 4969 2168 5021 2220
rect 5215 2168 5267 2220
rect 5543 2016 5595 2068
rect 5889 2016 5941 2068
rect 5461 1242 5513 1294
rect 5971 1242 6023 1294
rect 6217 2168 6269 2220
rect 1729 404 1781 456
rect 2215 404 2267 456
rect 2977 404 3029 456
rect 3463 404 3515 456
rect 4225 404 4277 456
rect 4711 404 4763 456
rect 5473 404 5525 456
rect 5959 404 6011 456
rect 1729 82 1781 134
rect 2215 82 2267 134
rect 2977 82 3029 134
rect 3463 82 3515 134
rect 4225 82 4277 134
rect 4711 82 4763 134
rect 5473 82 5525 134
rect 5959 82 6011 134
<< metal2 >>
rect 1469 2222 1525 2231
rect 1469 2157 1525 2166
rect 2471 2222 2527 2231
rect 2471 2157 2527 2166
rect 2717 2222 2773 2231
rect 2717 2157 2773 2166
rect 3719 2222 3775 2231
rect 3719 2157 3775 2166
rect 3965 2222 4021 2231
rect 3965 2157 4021 2166
rect 4967 2222 5023 2231
rect 4967 2157 5023 2166
rect 5213 2222 5269 2231
rect 5213 2157 5269 2166
rect 6215 2222 6271 2231
rect 6215 2157 6271 2166
rect 1797 2070 1853 2079
rect 1797 2005 1853 2014
rect 2143 2070 2199 2079
rect 2143 2005 2199 2014
rect 3045 2070 3101 2079
rect 3045 2005 3101 2014
rect 3391 2070 3447 2079
rect 3391 2005 3447 2014
rect 4293 2070 4349 2079
rect 4293 2005 4349 2014
rect 4639 2070 4695 2079
rect 4639 2005 4695 2014
rect 5541 2070 5597 2079
rect 5541 2005 5597 2014
rect 5887 2070 5943 2079
rect 5887 2005 5943 2014
rect 1715 1296 1771 1305
rect 1715 1231 1771 1240
rect 2225 1296 2281 1305
rect 2225 1231 2281 1240
rect 2963 1296 3019 1305
rect 2963 1231 3019 1240
rect 3473 1296 3529 1305
rect 3473 1231 3529 1240
rect 4211 1296 4267 1305
rect 4211 1231 4267 1240
rect 4721 1296 4777 1305
rect 4721 1231 4777 1240
rect 5459 1296 5515 1305
rect 5459 1231 5515 1240
rect 5969 1296 6025 1305
rect 5969 1231 6025 1240
rect 1727 458 1783 467
rect 1727 393 1783 402
rect 2213 458 2269 467
rect 2213 393 2269 402
rect 2975 458 3031 467
rect 2975 393 3031 402
rect 3461 458 3517 467
rect 3461 393 3517 402
rect 4223 458 4279 467
rect 4223 393 4279 402
rect 4709 458 4765 467
rect 4709 393 4765 402
rect 5471 458 5527 467
rect 5471 393 5527 402
rect 5957 458 6013 467
rect 5957 393 6013 402
rect 1727 136 1783 145
rect 1727 71 1783 80
rect 2213 136 2269 145
rect 2213 71 2269 80
rect 2975 136 3031 145
rect 2975 71 3031 80
rect 3461 136 3517 145
rect 3461 71 3517 80
rect 4223 136 4279 145
rect 4223 71 4279 80
rect 4709 136 4765 145
rect 4709 71 4765 80
rect 5471 136 5527 145
rect 5471 71 5527 80
rect 5957 136 6013 145
rect 5957 71 6013 80
<< via2 >>
rect 1469 2220 1525 2222
rect 1469 2168 1471 2220
rect 1471 2168 1523 2220
rect 1523 2168 1525 2220
rect 1469 2166 1525 2168
rect 2471 2220 2527 2222
rect 2471 2168 2473 2220
rect 2473 2168 2525 2220
rect 2525 2168 2527 2220
rect 2471 2166 2527 2168
rect 2717 2220 2773 2222
rect 2717 2168 2719 2220
rect 2719 2168 2771 2220
rect 2771 2168 2773 2220
rect 2717 2166 2773 2168
rect 3719 2220 3775 2222
rect 3719 2168 3721 2220
rect 3721 2168 3773 2220
rect 3773 2168 3775 2220
rect 3719 2166 3775 2168
rect 3965 2220 4021 2222
rect 3965 2168 3967 2220
rect 3967 2168 4019 2220
rect 4019 2168 4021 2220
rect 3965 2166 4021 2168
rect 4967 2220 5023 2222
rect 4967 2168 4969 2220
rect 4969 2168 5021 2220
rect 5021 2168 5023 2220
rect 4967 2166 5023 2168
rect 5213 2220 5269 2222
rect 5213 2168 5215 2220
rect 5215 2168 5267 2220
rect 5267 2168 5269 2220
rect 5213 2166 5269 2168
rect 6215 2220 6271 2222
rect 6215 2168 6217 2220
rect 6217 2168 6269 2220
rect 6269 2168 6271 2220
rect 6215 2166 6271 2168
rect 1797 2068 1853 2070
rect 1797 2016 1799 2068
rect 1799 2016 1851 2068
rect 1851 2016 1853 2068
rect 1797 2014 1853 2016
rect 2143 2068 2199 2070
rect 2143 2016 2145 2068
rect 2145 2016 2197 2068
rect 2197 2016 2199 2068
rect 2143 2014 2199 2016
rect 3045 2068 3101 2070
rect 3045 2016 3047 2068
rect 3047 2016 3099 2068
rect 3099 2016 3101 2068
rect 3045 2014 3101 2016
rect 3391 2068 3447 2070
rect 3391 2016 3393 2068
rect 3393 2016 3445 2068
rect 3445 2016 3447 2068
rect 3391 2014 3447 2016
rect 4293 2068 4349 2070
rect 4293 2016 4295 2068
rect 4295 2016 4347 2068
rect 4347 2016 4349 2068
rect 4293 2014 4349 2016
rect 4639 2068 4695 2070
rect 4639 2016 4641 2068
rect 4641 2016 4693 2068
rect 4693 2016 4695 2068
rect 4639 2014 4695 2016
rect 5541 2068 5597 2070
rect 5541 2016 5543 2068
rect 5543 2016 5595 2068
rect 5595 2016 5597 2068
rect 5541 2014 5597 2016
rect 5887 2068 5943 2070
rect 5887 2016 5889 2068
rect 5889 2016 5941 2068
rect 5941 2016 5943 2068
rect 5887 2014 5943 2016
rect 1715 1294 1771 1296
rect 1715 1242 1717 1294
rect 1717 1242 1769 1294
rect 1769 1242 1771 1294
rect 1715 1240 1771 1242
rect 2225 1294 2281 1296
rect 2225 1242 2227 1294
rect 2227 1242 2279 1294
rect 2279 1242 2281 1294
rect 2225 1240 2281 1242
rect 2963 1294 3019 1296
rect 2963 1242 2965 1294
rect 2965 1242 3017 1294
rect 3017 1242 3019 1294
rect 2963 1240 3019 1242
rect 3473 1294 3529 1296
rect 3473 1242 3475 1294
rect 3475 1242 3527 1294
rect 3527 1242 3529 1294
rect 3473 1240 3529 1242
rect 4211 1294 4267 1296
rect 4211 1242 4213 1294
rect 4213 1242 4265 1294
rect 4265 1242 4267 1294
rect 4211 1240 4267 1242
rect 4721 1294 4777 1296
rect 4721 1242 4723 1294
rect 4723 1242 4775 1294
rect 4775 1242 4777 1294
rect 4721 1240 4777 1242
rect 5459 1294 5515 1296
rect 5459 1242 5461 1294
rect 5461 1242 5513 1294
rect 5513 1242 5515 1294
rect 5459 1240 5515 1242
rect 5969 1294 6025 1296
rect 5969 1242 5971 1294
rect 5971 1242 6023 1294
rect 6023 1242 6025 1294
rect 5969 1240 6025 1242
rect 1727 456 1783 458
rect 1727 404 1729 456
rect 1729 404 1781 456
rect 1781 404 1783 456
rect 1727 402 1783 404
rect 2213 456 2269 458
rect 2213 404 2215 456
rect 2215 404 2267 456
rect 2267 404 2269 456
rect 2213 402 2269 404
rect 2975 456 3031 458
rect 2975 404 2977 456
rect 2977 404 3029 456
rect 3029 404 3031 456
rect 2975 402 3031 404
rect 3461 456 3517 458
rect 3461 404 3463 456
rect 3463 404 3515 456
rect 3515 404 3517 456
rect 3461 402 3517 404
rect 4223 456 4279 458
rect 4223 404 4225 456
rect 4225 404 4277 456
rect 4277 404 4279 456
rect 4223 402 4279 404
rect 4709 456 4765 458
rect 4709 404 4711 456
rect 4711 404 4763 456
rect 4763 404 4765 456
rect 4709 402 4765 404
rect 5471 456 5527 458
rect 5471 404 5473 456
rect 5473 404 5525 456
rect 5525 404 5527 456
rect 5471 402 5527 404
rect 5957 456 6013 458
rect 5957 404 5959 456
rect 5959 404 6011 456
rect 6011 404 6013 456
rect 5957 402 6013 404
rect 1727 134 1783 136
rect 1727 82 1729 134
rect 1729 82 1781 134
rect 1781 82 1783 134
rect 1727 80 1783 82
rect 2213 134 2269 136
rect 2213 82 2215 134
rect 2215 82 2267 134
rect 2267 82 2269 134
rect 2213 80 2269 82
rect 2975 134 3031 136
rect 2975 82 2977 134
rect 2977 82 3029 134
rect 3029 82 3031 134
rect 2975 80 3031 82
rect 3461 134 3517 136
rect 3461 82 3463 134
rect 3463 82 3515 134
rect 3515 82 3517 134
rect 3461 80 3517 82
rect 4223 134 4279 136
rect 4223 82 4225 134
rect 4225 82 4277 134
rect 4277 82 4279 134
rect 4223 80 4279 82
rect 4709 134 4765 136
rect 4709 82 4711 134
rect 4711 82 4763 134
rect 4763 82 4765 134
rect 4709 80 4765 82
rect 5471 134 5527 136
rect 5471 82 5473 134
rect 5473 82 5525 134
rect 5525 82 5527 134
rect 5471 80 5527 82
rect 5957 134 6013 136
rect 5957 82 5959 134
rect 5959 82 6011 134
rect 6011 82 6013 134
rect 5957 80 6013 82
<< metal3 >>
rect 1464 2224 1530 2227
rect 2466 2224 2532 2227
rect 2712 2224 2778 2227
rect 3714 2224 3780 2227
rect 3960 2224 4026 2227
rect 4962 2224 5028 2227
rect 5208 2224 5274 2227
rect 6210 2224 6276 2227
rect 0 2222 6366 2224
rect 0 2166 1469 2222
rect 1525 2166 2471 2222
rect 2527 2166 2717 2222
rect 2773 2166 3719 2222
rect 3775 2166 3965 2222
rect 4021 2166 4967 2222
rect 5023 2166 5213 2222
rect 5269 2166 6215 2222
rect 6271 2166 6366 2222
rect 0 2164 6366 2166
rect 1464 2161 1530 2164
rect 2466 2161 2532 2164
rect 2712 2161 2778 2164
rect 3714 2161 3780 2164
rect 3960 2161 4026 2164
rect 4962 2161 5028 2164
rect 5208 2161 5274 2164
rect 6210 2161 6276 2164
rect 1776 2070 1874 2091
rect 1776 2014 1797 2070
rect 1853 2014 1874 2070
rect 1776 1993 1874 2014
rect 2122 2070 2220 2091
rect 2122 2014 2143 2070
rect 2199 2014 2220 2070
rect 2122 1993 2220 2014
rect 3024 2070 3122 2091
rect 3024 2014 3045 2070
rect 3101 2014 3122 2070
rect 3024 1993 3122 2014
rect 3370 2070 3468 2091
rect 3370 2014 3391 2070
rect 3447 2014 3468 2070
rect 3370 1993 3468 2014
rect 4272 2070 4370 2091
rect 4272 2014 4293 2070
rect 4349 2014 4370 2070
rect 4272 1993 4370 2014
rect 4618 2070 4716 2091
rect 4618 2014 4639 2070
rect 4695 2014 4716 2070
rect 4618 1993 4716 2014
rect 5520 2070 5618 2091
rect 5520 2014 5541 2070
rect 5597 2014 5618 2070
rect 5520 1993 5618 2014
rect 5866 2070 5964 2091
rect 5866 2014 5887 2070
rect 5943 2014 5964 2070
rect 5866 1993 5964 2014
rect 1694 1296 1792 1317
rect 1694 1240 1715 1296
rect 1771 1240 1792 1296
rect 1694 1219 1792 1240
rect 2204 1296 2302 1317
rect 2204 1240 2225 1296
rect 2281 1240 2302 1296
rect 2204 1219 2302 1240
rect 2942 1296 3040 1317
rect 2942 1240 2963 1296
rect 3019 1240 3040 1296
rect 2942 1219 3040 1240
rect 3452 1296 3550 1317
rect 3452 1240 3473 1296
rect 3529 1240 3550 1296
rect 3452 1219 3550 1240
rect 4190 1296 4288 1317
rect 4190 1240 4211 1296
rect 4267 1240 4288 1296
rect 4190 1219 4288 1240
rect 4700 1296 4798 1317
rect 4700 1240 4721 1296
rect 4777 1240 4798 1296
rect 4700 1219 4798 1240
rect 5438 1296 5536 1317
rect 5438 1240 5459 1296
rect 5515 1240 5536 1296
rect 5438 1219 5536 1240
rect 5948 1296 6046 1317
rect 5948 1240 5969 1296
rect 6025 1240 6046 1296
rect 5948 1219 6046 1240
rect 1706 458 1804 479
rect 1706 402 1727 458
rect 1783 402 1804 458
rect 1706 381 1804 402
rect 2192 458 2290 479
rect 2192 402 2213 458
rect 2269 402 2290 458
rect 2192 381 2290 402
rect 2954 458 3052 479
rect 2954 402 2975 458
rect 3031 402 3052 458
rect 2954 381 3052 402
rect 3440 458 3538 479
rect 3440 402 3461 458
rect 3517 402 3538 458
rect 3440 381 3538 402
rect 4202 458 4300 479
rect 4202 402 4223 458
rect 4279 402 4300 458
rect 4202 381 4300 402
rect 4688 458 4786 479
rect 4688 402 4709 458
rect 4765 402 4786 458
rect 4688 381 4786 402
rect 5450 458 5548 479
rect 5450 402 5471 458
rect 5527 402 5548 458
rect 5450 381 5548 402
rect 5936 458 6034 479
rect 5936 402 5957 458
rect 6013 402 6034 458
rect 5936 381 6034 402
rect 1706 136 1804 157
rect 1706 80 1727 136
rect 1783 80 1804 136
rect 1706 59 1804 80
rect 2192 136 2290 157
rect 2192 80 2213 136
rect 2269 80 2290 136
rect 2192 59 2290 80
rect 2954 136 3052 157
rect 2954 80 2975 136
rect 3031 80 3052 136
rect 2954 59 3052 80
rect 3440 136 3538 157
rect 3440 80 3461 136
rect 3517 80 3538 136
rect 3440 59 3538 80
rect 4202 136 4300 157
rect 4202 80 4223 136
rect 4279 80 4300 136
rect 4202 59 4300 80
rect 4688 136 4786 157
rect 4688 80 4709 136
rect 4765 80 4786 136
rect 4688 59 4786 80
rect 5450 136 5548 157
rect 5450 80 5471 136
rect 5527 80 5548 136
rect 5450 59 5548 80
rect 5936 136 6034 157
rect 5936 80 5957 136
rect 6013 80 6034 136
rect 5936 59 6034 80
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 6210 0 1 2157
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 6211 0 1 2162
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 5208 0 1 2157
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 5209 0 1 2162
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 4962 0 1 2157
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 4963 0 1 2162
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 3960 0 1 2157
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 3961 0 1 2162
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 3714 0 1 2157
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 3715 0 1 2162
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 2712 0 1 2157
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 2713 0 1 2162
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 2466 0 1 2157
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 2467 0 1 2162
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 1464 0 1 2157
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 1465 0 1 2162
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 5952 0 1 393
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 5953 0 1 398
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 5964 0 1 1231
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 5965 0 1 1236
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 5952 0 1 71
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 5953 0 1 76
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 5882 0 1 2005
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 5883 0 1 2010
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 5466 0 1 393
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 5467 0 1 398
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 5454 0 1 1231
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 5455 0 1 1236
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 5466 0 1 71
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 5467 0 1 76
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 5536 0 1 2005
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 5537 0 1 2010
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 4704 0 1 393
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1634918361
transform 1 0 4705 0 1 398
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1634918361
transform 1 0 4716 0 1 1231
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1634918361
transform 1 0 4717 0 1 1236
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1634918361
transform 1 0 4704 0 1 71
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1634918361
transform 1 0 4705 0 1 76
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1634918361
transform 1 0 4634 0 1 2005
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1634918361
transform 1 0 4635 0 1 2010
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1634918361
transform 1 0 4218 0 1 393
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1634918361
transform 1 0 4219 0 1 398
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1634918361
transform 1 0 4206 0 1 1231
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1634918361
transform 1 0 4207 0 1 1236
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1634918361
transform 1 0 4218 0 1 71
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1634918361
transform 1 0 4219 0 1 76
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1634918361
transform 1 0 4288 0 1 2005
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1634918361
transform 1 0 4289 0 1 2010
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1634918361
transform 1 0 3456 0 1 393
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1634918361
transform 1 0 3457 0 1 398
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1634918361
transform 1 0 3468 0 1 1231
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1634918361
transform 1 0 3469 0 1 1236
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1634918361
transform 1 0 3456 0 1 71
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1634918361
transform 1 0 3457 0 1 76
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1634918361
transform 1 0 3386 0 1 2005
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1634918361
transform 1 0 3387 0 1 2010
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1634918361
transform 1 0 2970 0 1 393
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1634918361
transform 1 0 2971 0 1 398
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1634918361
transform 1 0 2958 0 1 1231
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1634918361
transform 1 0 2959 0 1 1236
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1634918361
transform 1 0 2970 0 1 71
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1634918361
transform 1 0 2971 0 1 76
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1634918361
transform 1 0 3040 0 1 2005
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1634918361
transform 1 0 3041 0 1 2010
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1634918361
transform 1 0 2208 0 1 393
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1634918361
transform 1 0 2209 0 1 398
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1634918361
transform 1 0 2220 0 1 1231
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1634918361
transform 1 0 2221 0 1 1236
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1634918361
transform 1 0 2208 0 1 71
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1634918361
transform 1 0 2209 0 1 76
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1634918361
transform 1 0 2138 0 1 2005
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1634918361
transform 1 0 2139 0 1 2010
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1634918361
transform 1 0 1722 0 1 393
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1634918361
transform 1 0 1723 0 1 398
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1634918361
transform 1 0 1710 0 1 1231
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1634918361
transform 1 0 1711 0 1 1236
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1634918361
transform 1 0 1722 0 1 71
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1634918361
transform 1 0 1723 0 1 76
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1634918361
transform 1 0 1792 0 1 2005
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1634918361
transform 1 0 1793 0 1 2010
box 0 0 1 1
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_0
timestamp 1634918361
transform -1 0 6366 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_1
timestamp 1634918361
transform 1 0 5118 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_2
timestamp 1634918361
transform -1 0 5118 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_3
timestamp 1634918361
transform 1 0 3870 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_4
timestamp 1634918361
transform -1 0 3870 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_5
timestamp 1634918361
transform 1 0 2622 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_6
timestamp 1634918361
transform -1 0 2622 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_7
timestamp 1634918361
transform 1 0 1374 0 1 0
box -541 0 937 2256
<< labels >>
rlabel metal3 s 2122 1993 2220 2091 4 gnd
port 1 nsew
rlabel metal3 s 5866 1993 5964 2091 4 gnd
port 1 nsew
rlabel metal3 s 3440 59 3538 157 4 gnd
port 1 nsew
rlabel metal3 s 3370 1993 3468 2091 4 gnd
port 1 nsew
rlabel metal3 s 5936 59 6034 157 4 gnd
port 1 nsew
rlabel metal3 s 5520 1993 5618 2091 4 gnd
port 1 nsew
rlabel metal3 s 5450 59 5548 157 4 gnd
port 1 nsew
rlabel metal3 s 4272 1993 4370 2091 4 gnd
port 1 nsew
rlabel metal3 s 2954 59 3052 157 4 gnd
port 1 nsew
rlabel metal3 s 4202 59 4300 157 4 gnd
port 1 nsew
rlabel metal3 s 4618 1993 4716 2091 4 gnd
port 1 nsew
rlabel metal3 s 1706 59 1804 157 4 gnd
port 1 nsew
rlabel metal3 s 4688 59 4786 157 4 gnd
port 1 nsew
rlabel metal3 s 2192 59 2290 157 4 gnd
port 1 nsew
rlabel metal3 s 1776 1993 1874 2091 4 gnd
port 1 nsew
rlabel metal3 s 3024 1993 3122 2091 4 gnd
port 1 nsew
rlabel metal3 s 3452 1219 3550 1317 4 vdd
port 2 nsew
rlabel metal3 s 2942 1219 3040 1317 4 vdd
port 2 nsew
rlabel metal3 s 1706 381 1804 479 4 vdd
port 2 nsew
rlabel metal3 s 4700 1219 4798 1317 4 vdd
port 2 nsew
rlabel metal3 s 3440 381 3538 479 4 vdd
port 2 nsew
rlabel metal3 s 4202 381 4300 479 4 vdd
port 2 nsew
rlabel metal3 s 5936 381 6034 479 4 vdd
port 2 nsew
rlabel metal3 s 5948 1219 6046 1317 4 vdd
port 2 nsew
rlabel metal3 s 5450 381 5548 479 4 vdd
port 2 nsew
rlabel metal3 s 2192 381 2290 479 4 vdd
port 2 nsew
rlabel metal3 s 4190 1219 4288 1317 4 vdd
port 2 nsew
rlabel metal3 s 4688 381 4786 479 4 vdd
port 2 nsew
rlabel metal3 s 1694 1219 1792 1317 4 vdd
port 2 nsew
rlabel metal3 s 2954 381 3052 479 4 vdd
port 2 nsew
rlabel metal3 s 2204 1219 2302 1317 4 vdd
port 2 nsew
rlabel metal3 s 5438 1219 5536 1317 4 vdd
port 2 nsew
rlabel metal1 s 1570 1130 1604 2256 4 bl_0
port 3 nsew
rlabel metal1 s 1646 1142 1674 2256 4 br_0
port 4 nsew
rlabel metal1 s 1478 0 1524 254 4 data_0
port 5 nsew
rlabel metal1 s 2392 1130 2426 2256 4 bl_1
port 6 nsew
rlabel metal1 s 2322 1142 2350 2256 4 br_1
port 7 nsew
rlabel metal1 s 2472 0 2518 254 4 data_1
port 8 nsew
rlabel metal1 s 2818 1130 2852 2256 4 bl_2
port 9 nsew
rlabel metal1 s 2894 1142 2922 2256 4 br_2
port 10 nsew
rlabel metal1 s 2726 0 2772 254 4 data_2
port 11 nsew
rlabel metal1 s 3640 1130 3674 2256 4 bl_3
port 12 nsew
rlabel metal1 s 3570 1142 3598 2256 4 br_3
port 13 nsew
rlabel metal1 s 3720 0 3766 254 4 data_3
port 14 nsew
rlabel metal1 s 4066 1130 4100 2256 4 bl_4
port 15 nsew
rlabel metal1 s 4142 1142 4170 2256 4 br_4
port 16 nsew
rlabel metal1 s 3974 0 4020 254 4 data_4
port 17 nsew
rlabel metal1 s 4888 1130 4922 2256 4 bl_5
port 18 nsew
rlabel metal1 s 4818 1142 4846 2256 4 br_5
port 19 nsew
rlabel metal1 s 4968 0 5014 254 4 data_5
port 20 nsew
rlabel metal1 s 5314 1130 5348 2256 4 bl_6
port 21 nsew
rlabel metal1 s 5390 1142 5418 2256 4 br_6
port 22 nsew
rlabel metal1 s 5222 0 5268 254 4 data_6
port 23 nsew
rlabel metal1 s 6136 1130 6170 2256 4 bl_7
port 24 nsew
rlabel metal1 s 6066 1142 6094 2256 4 br_7
port 25 nsew
rlabel metal1 s 6216 0 6262 254 4 data_7
port 26 nsew
rlabel metal3 s 0 2164 6366 2224 4 en
port 27 nsew
<< properties >>
string FIXED_BBOX 0 0 6366 2256
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 824536
string GDS_START 808136
<< end >>
