magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1190 -1316 2896 1750
<< locali >>
rect 70 282 136 316
rect 549 314 970 348
rect 70 174 136 208
rect 936 170 970 314
rect 1041 103 1618 137
<< metal1 >>
rect 246 -30 294 402
rect 670 -32 720 402
rect 1060 0 1088 395
rect 1456 0 1484 395
use pinv_dec  pinv_dec_0
timestamp 1634918361
transform 1 0 876 0 1 0
box 44 0 760 490
use sky130_fd_bd_sram__openram_dp_nand2_dec  sky130_fd_bd_sram__openram_dp_nand2_dec_0
timestamp 1634918361
transform 1 0 0 0 1 0
box 70 -56 888 476
<< labels >>
rlabel locali s 1329 120 1329 120 4 Z
port 1 nsew
rlabel locali s 103 299 103 299 4 A
port 2 nsew
rlabel locali s 103 191 103 191 4 B
port 3 nsew
rlabel metal1 s 1456 0 1484 395 4 vdd
port 4 nsew
rlabel metal1 s 670 -32 720 402 4 vdd
port 4 nsew
rlabel metal1 s 246 -30 294 402 4 gnd
port 5 nsew
rlabel metal1 s 1060 0 1088 395 4 gnd
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1618 395
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 986614
string GDS_START 985162
<< end >>
