magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1309 -1022 8167 8458
<< locali >>
rect 1931 6644 1965 6660
rect 1931 6594 1965 6610
rect 3179 6644 3213 6660
rect 3179 6594 3213 6610
rect 4427 6644 4461 6660
rect 4427 6594 4461 6610
rect 5675 6644 5709 6660
rect 5675 6594 5709 6610
<< viali >>
rect 1931 6610 1965 6644
rect 3179 6610 3213 6644
rect 4427 6610 4461 6644
rect 5675 6610 5709 6644
<< metal1 >>
rect 1919 6644 1977 6650
rect 1919 6610 1931 6644
rect 1965 6641 1977 6644
rect 2382 6641 2388 6653
rect 1965 6613 2388 6641
rect 1965 6610 1977 6613
rect 1919 6604 1977 6610
rect 2382 6601 2388 6613
rect 2440 6601 2446 6653
rect 3167 6644 3225 6650
rect 3167 6610 3179 6644
rect 3213 6641 3225 6644
rect 3630 6641 3636 6653
rect 3213 6613 3636 6641
rect 3213 6610 3225 6613
rect 3167 6604 3225 6610
rect 3630 6601 3636 6613
rect 3688 6601 3694 6653
rect 4415 6644 4473 6650
rect 4415 6610 4427 6644
rect 4461 6641 4473 6644
rect 4878 6641 4884 6653
rect 4461 6613 4884 6641
rect 4461 6610 4473 6613
rect 4415 6604 4473 6610
rect 4878 6601 4884 6613
rect 4936 6601 4942 6653
rect 5663 6644 5721 6650
rect 5663 6610 5675 6644
rect 5709 6641 5721 6644
rect 6126 6641 6132 6653
rect 5709 6613 6132 6641
rect 5709 6610 5721 6613
rect 5663 6604 5721 6610
rect 6126 6601 6132 6613
rect 6184 6601 6190 6653
rect 1629 5717 1689 5773
rect 2183 5717 2243 5773
rect 2877 5717 2937 5773
rect 3431 5717 3491 5773
rect 4125 5717 4185 5773
rect 4679 5717 4739 5773
rect 5373 5717 5433 5773
rect 5927 5717 5987 5773
rect 2382 5683 2388 5692
rect 1473 5649 2388 5683
rect 2382 5640 2388 5649
rect 2440 5683 2446 5692
rect 3630 5683 3636 5692
rect 2440 5649 2498 5683
rect 2721 5649 3636 5683
rect 2440 5640 2446 5649
rect 3630 5640 3636 5649
rect 3688 5683 3694 5692
rect 4878 5683 4884 5692
rect 3688 5649 3746 5683
rect 3969 5649 4884 5683
rect 3688 5640 3694 5649
rect 4878 5640 4884 5649
rect 4936 5683 4942 5692
rect 6126 5683 6132 5692
rect 4936 5649 4994 5683
rect 5217 5649 6132 5683
rect 4936 5640 4942 5649
rect 6126 5640 6132 5649
rect 6184 5683 6190 5692
rect 6184 5649 6242 5683
rect 6184 5640 6190 5649
rect 1501 3700 1529 3766
rect 1501 3672 1601 3700
rect 1478 3260 1524 3514
rect 1573 2384 1601 3672
rect 1703 3620 1731 3766
rect 1646 3592 1731 3620
rect 2141 3620 2169 3766
rect 2343 3700 2371 3766
rect 2749 3700 2777 3766
rect 2343 3672 2423 3700
rect 2749 3672 2849 3700
rect 2141 3592 2350 3620
rect 1646 2372 1674 3592
rect 2322 2372 2350 3592
rect 2395 2384 2423 3672
rect 2472 3260 2518 3514
rect 2726 3260 2772 3514
rect 2821 2384 2849 3672
rect 2951 3620 2979 3766
rect 2894 3592 2979 3620
rect 3389 3620 3417 3766
rect 3591 3700 3619 3766
rect 3997 3700 4025 3766
rect 3591 3672 3671 3700
rect 3997 3672 4097 3700
rect 3389 3592 3598 3620
rect 2894 2372 2922 3592
rect 3570 2372 3598 3592
rect 3643 2384 3671 3672
rect 3720 3260 3766 3514
rect 3974 3260 4020 3514
rect 4069 2384 4097 3672
rect 4199 3620 4227 3766
rect 4142 3592 4227 3620
rect 4637 3620 4665 3766
rect 4839 3700 4867 3766
rect 5245 3700 5273 3766
rect 4839 3672 4919 3700
rect 5245 3672 5345 3700
rect 4637 3592 4846 3620
rect 4142 2372 4170 3592
rect 4818 2372 4846 3592
rect 4891 2384 4919 3672
rect 4968 3260 5014 3514
rect 5222 3260 5268 3514
rect 5317 2384 5345 3672
rect 5447 3620 5475 3766
rect 5390 3592 5475 3620
rect 5885 3620 5913 3766
rect 6087 3700 6115 3766
rect 6087 3672 6167 3700
rect 5885 3592 6094 3620
rect 5390 2372 5418 3592
rect 6066 2372 6094 3592
rect 6139 2384 6167 3672
rect 6216 3260 6262 3514
rect 1573 1192 1601 1258
rect 1440 1164 1601 1192
rect 816 252 844 1006
rect 1280 252 1308 1006
rect 1440 252 1468 1164
rect 1646 1112 1674 1258
rect 2322 1112 2350 1258
rect 2395 1192 2423 1258
rect 2821 1192 2849 1258
rect 2395 1164 2556 1192
rect 1646 1084 1932 1112
rect 1904 252 1932 1084
rect 2064 1084 2350 1112
rect 2064 252 2092 1084
rect 2528 252 2556 1164
rect 2688 1164 2849 1192
rect 2688 252 2716 1164
rect 2894 1112 2922 1258
rect 3570 1112 3598 1258
rect 3643 1192 3671 1258
rect 4069 1192 4097 1258
rect 3643 1164 3804 1192
rect 2894 1084 3180 1112
rect 3152 252 3180 1084
rect 3312 1084 3598 1112
rect 3312 252 3340 1084
rect 3776 252 3804 1164
rect 3936 1164 4097 1192
rect 3936 252 3964 1164
rect 4142 1112 4170 1258
rect 4818 1112 4846 1258
rect 4891 1192 4919 1258
rect 5317 1192 5345 1258
rect 4891 1164 5052 1192
rect 4142 1084 4428 1112
rect 4400 252 4428 1084
rect 4560 1084 4846 1112
rect 4560 252 4588 1084
rect 5024 252 5052 1164
rect 5184 1164 5345 1192
rect 5184 252 5212 1164
rect 5390 1112 5418 1258
rect 6066 1112 6094 1258
rect 6139 1192 6167 1258
rect 6139 1164 6300 1192
rect 5390 1084 5676 1112
rect 5648 252 5676 1084
rect 5808 1084 6094 1112
rect 5808 252 5836 1084
rect 6272 252 6300 1164
<< via1 >>
rect 2388 6601 2440 6653
rect 3636 6601 3688 6653
rect 4884 6601 4936 6653
rect 6132 6601 6184 6653
rect 2388 5640 2440 5692
rect 3636 5640 3688 5692
rect 4884 5640 4936 5692
rect 6132 5640 6184 5692
<< metal2 >>
rect 1360 6865 1388 6893
rect 2608 6865 2636 6893
rect 3856 6865 3884 6893
rect 5104 6865 5132 6893
rect 2388 6653 2440 6659
rect 2388 6595 2440 6601
rect 3636 6653 3688 6659
rect 3636 6595 3688 6601
rect 4884 6653 4936 6659
rect 4884 6595 4936 6601
rect 6132 6653 6184 6659
rect 6132 6595 6184 6601
rect 2400 5698 2428 6595
rect 3648 5698 3676 6595
rect 4896 5698 4924 6595
rect 6144 5698 6172 6595
rect 2388 5692 2440 5698
rect 2388 5634 2440 5640
rect 3636 5692 3688 5698
rect 3636 5634 3688 5640
rect 4884 5692 4936 5698
rect 4884 5634 4936 5640
rect 6132 5692 6184 5698
rect 6132 5634 6184 5640
<< metal3 >>
rect -49 7100 49 7198
rect 6317 7100 6415 7198
rect 0 6601 6366 6661
rect -49 5980 49 6078
rect 6317 5980 6415 6078
rect 1601 5537 1699 5635
rect 2173 5537 2271 5635
rect 2849 5537 2947 5635
rect 3421 5537 3519 5635
rect 4097 5537 4195 5635
rect 4669 5537 4767 5635
rect 5345 5537 5443 5635
rect 5917 5537 6015 5635
rect 1587 5121 1685 5219
rect 2187 5121 2285 5219
rect 2835 5121 2933 5219
rect 3435 5121 3533 5219
rect 4083 5121 4181 5219
rect 4683 5121 4781 5219
rect 5331 5121 5429 5219
rect 5931 5121 6029 5219
rect 1702 4919 1800 5017
rect 2072 4919 2170 5017
rect 2950 4919 3048 5017
rect 3320 4919 3418 5017
rect 4198 4919 4296 5017
rect 4568 4919 4666 5017
rect 5446 4919 5544 5017
rect 5816 4919 5914 5017
rect 1581 4587 1679 4685
rect 2193 4587 2291 4685
rect 2829 4587 2927 4685
rect 3441 4587 3539 4685
rect 4077 4587 4175 4685
rect 4689 4587 4787 4685
rect 5325 4587 5423 4685
rect 5937 4587 6035 4685
rect 1592 4150 1690 4248
rect 2182 4150 2280 4248
rect 2840 4150 2938 4248
rect 3430 4150 3528 4248
rect 4088 4150 4186 4248
rect 4678 4150 4776 4248
rect 5336 4150 5434 4248
rect 5926 4150 6024 4248
rect 1706 3357 1804 3455
rect 2192 3357 2290 3455
rect 2954 3357 3052 3455
rect 3440 3357 3538 3455
rect 4202 3357 4300 3455
rect 4688 3357 4786 3455
rect 5450 3357 5548 3455
rect 5936 3357 6034 3455
rect 1706 3035 1804 3133
rect 2192 3035 2290 3133
rect 2954 3035 3052 3133
rect 3440 3035 3538 3133
rect 4202 3035 4300 3133
rect 4688 3035 4786 3133
rect 5450 3035 5548 3133
rect 5936 3035 6034 3133
rect 1694 2197 1792 2295
rect 2204 2197 2302 2295
rect 2942 2197 3040 2295
rect 3452 2197 3550 2295
rect 4190 2197 4288 2295
rect 4700 2197 4798 2295
rect 5438 2197 5536 2295
rect 5948 2197 6046 2295
rect 1776 1423 1874 1521
rect 2122 1423 2220 1521
rect 3024 1423 3122 1521
rect 3370 1423 3468 1521
rect 4272 1423 4370 1521
rect 4618 1423 4716 1521
rect 5520 1423 5618 1521
rect 5866 1423 5964 1521
rect 0 1290 6366 1350
rect 0 951 6366 1011
rect 1132 313 1230 411
rect 1518 313 1616 411
rect 2380 313 2478 411
rect 2766 313 2864 411
rect 3628 313 3726 411
rect 4014 313 4112 411
rect 4876 313 4974 411
rect 5262 313 5360 411
rect 6124 313 6222 411
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 6126 0 1 6595
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 6126 0 1 5634
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 5663 0 1 6594
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 4878 0 1 6595
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 4878 0 1 5634
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 4415 0 1 6594
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 3630 0 1 6595
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 3630 0 1 5634
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 3167 0 1 6594
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 2382 0 1 6595
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 2382 0 1 5634
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 1919 0 1 6594
box 0 0 1 1
use write_mask_and_array  write_mask_and_array_0
timestamp 1634918361
transform 1 0 0 0 -1 7149
box -49 -49 6415 1177
use write_driver_array  write_driver_array_0
timestamp 1634918361
transform 1 0 0 0 -1 5777
box 998 4 6618 2011
use sense_amp_array  sense_amp_array_0
timestamp 1634918361
transform 1 0 0 0 -1 3514
box 0 0 6907 2256
use precharge_array  precharge_array_0
timestamp 1634918361
transform 1 0 0 0 -1 1006
box 0 -12 6366 768
<< labels >>
rlabel metal2 s 1360 6865 1388 6893 4 bank_wmask_0
port 1 nsew
rlabel metal2 s 2608 6865 2636 6893 4 bank_wmask_1
port 2 nsew
rlabel metal2 s 3856 6865 3884 6893 4 bank_wmask_2
port 3 nsew
rlabel metal2 s 5104 6865 5132 6893 4 bank_wmask_3
port 4 nsew
rlabel locali s 1948 6627 1948 6627 4 wdriver_sel_0
port 5 nsew
rlabel metal1 s 1473 5649 2498 5683 4 wdriver_sel_0
port 5 nsew
rlabel metal1 s 2721 5649 3746 5683 4 wdriver_sel_1
port 6 nsew
rlabel locali s 3196 6627 3196 6627 4 wdriver_sel_1
port 6 nsew
rlabel metal1 s 3969 5649 4994 5683 4 wdriver_sel_2
port 7 nsew
rlabel locali s 4444 6627 4444 6627 4 wdriver_sel_2
port 7 nsew
rlabel locali s 5692 6627 5692 6627 4 wdriver_sel_3
port 8 nsew
rlabel metal1 s 5217 5649 6242 5683 4 wdriver_sel_3
port 8 nsew
rlabel metal1 s 1629 5717 1689 5773 4 din_0
port 9 nsew
rlabel metal1 s 2183 5717 2243 5773 4 din_1
port 10 nsew
rlabel metal1 s 2877 5717 2937 5773 4 din_2
port 11 nsew
rlabel metal1 s 3431 5717 3491 5773 4 din_3
port 12 nsew
rlabel metal1 s 4125 5717 4185 5773 4 din_4
port 13 nsew
rlabel metal1 s 4679 5717 4739 5773 4 din_5
port 14 nsew
rlabel metal1 s 5373 5717 5433 5773 4 din_6
port 15 nsew
rlabel metal1 s 5927 5717 5987 5773 4 din_7
port 16 nsew
rlabel metal1 s 1478 3260 1524 3514 4 dout_0
port 17 nsew
rlabel metal1 s 2472 3260 2518 3514 4 dout_1
port 18 nsew
rlabel metal1 s 2726 3260 2772 3514 4 dout_2
port 19 nsew
rlabel metal1 s 3720 3260 3766 3514 4 dout_3
port 20 nsew
rlabel metal1 s 3974 3260 4020 3514 4 dout_4
port 21 nsew
rlabel metal1 s 4968 3260 5014 3514 4 dout_5
port 22 nsew
rlabel metal1 s 5222 3260 5268 3514 4 dout_6
port 23 nsew
rlabel metal1 s 6216 3260 6262 3514 4 dout_7
port 24 nsew
rlabel metal1 s 1280 252 1308 1006 4 rbl_bl
port 25 nsew
rlabel metal1 s 816 252 844 1006 4 rbl_br
port 26 nsew
rlabel metal1 s 1440 252 1468 1006 4 bl_0
port 27 nsew
rlabel metal1 s 1904 252 1932 1006 4 br_0
port 28 nsew
rlabel metal1 s 2528 252 2556 1006 4 bl_1
port 29 nsew
rlabel metal1 s 2064 252 2092 1006 4 br_1
port 30 nsew
rlabel metal1 s 2688 252 2716 1006 4 bl_2
port 31 nsew
rlabel metal1 s 3152 252 3180 1006 4 br_2
port 32 nsew
rlabel metal1 s 3776 252 3804 1006 4 bl_3
port 33 nsew
rlabel metal1 s 3312 252 3340 1006 4 br_3
port 34 nsew
rlabel metal1 s 3936 252 3964 1006 4 bl_4
port 35 nsew
rlabel metal1 s 4400 252 4428 1006 4 br_4
port 36 nsew
rlabel metal1 s 5024 252 5052 1006 4 bl_5
port 37 nsew
rlabel metal1 s 4560 252 4588 1006 4 br_5
port 38 nsew
rlabel metal1 s 5184 252 5212 1006 4 bl_6
port 39 nsew
rlabel metal1 s 5648 252 5676 1006 4 br_6
port 40 nsew
rlabel metal1 s 6272 252 6300 1006 4 bl_7
port 41 nsew
rlabel metal1 s 5808 252 5836 1006 4 br_7
port 42 nsew
rlabel metal3 s 0 951 6366 1011 4 p_en_bar
port 43 nsew
rlabel metal3 s 0 1290 6366 1350 4 s_en
port 44 nsew
rlabel metal3 s 0 6601 6366 6661 4 w_en
port 45 nsew
rlabel metal3 s 2954 3035 3052 3133 4 vdd
port 46 nsew
rlabel metal3 s 3441 4587 3539 4685 4 vdd
port 46 nsew
rlabel metal3 s 3628 313 3726 411 4 vdd
port 46 nsew
rlabel metal3 s 5450 3035 5548 3133 4 vdd
port 46 nsew
rlabel metal3 s 5937 4587 6035 4685 4 vdd
port 46 nsew
rlabel metal3 s 5948 2197 6046 2295 4 vdd
port 46 nsew
rlabel metal3 s 2380 313 2478 411 4 vdd
port 46 nsew
rlabel metal3 s 5917 5537 6015 5635 4 vdd
port 46 nsew
rlabel metal3 s 1518 313 1616 411 4 vdd
port 46 nsew
rlabel metal3 s 2192 3035 2290 3133 4 vdd
port 46 nsew
rlabel metal3 s 2204 2197 2302 2295 4 vdd
port 46 nsew
rlabel metal3 s 5262 313 5360 411 4 vdd
port 46 nsew
rlabel metal3 s 2829 4587 2927 4685 4 vdd
port 46 nsew
rlabel metal3 s 3452 2197 3550 2295 4 vdd
port 46 nsew
rlabel metal3 s 4014 313 4112 411 4 vdd
port 46 nsew
rlabel metal3 s 3440 3035 3538 3133 4 vdd
port 46 nsew
rlabel metal3 s 5345 5537 5443 5635 4 vdd
port 46 nsew
rlabel metal3 s 4876 313 4974 411 4 vdd
port 46 nsew
rlabel metal3 s 1132 313 1230 411 4 vdd
port 46 nsew
rlabel metal3 s 4700 2197 4798 2295 4 vdd
port 46 nsew
rlabel metal3 s 2942 2197 3040 2295 4 vdd
port 46 nsew
rlabel metal3 s 4669 5537 4767 5635 4 vdd
port 46 nsew
rlabel metal3 s 4077 4587 4175 4685 4 vdd
port 46 nsew
rlabel metal3 s 2849 5537 2947 5635 4 vdd
port 46 nsew
rlabel metal3 s -49 5980 49 6078 4 vdd
port 46 nsew
rlabel metal3 s 5325 4587 5423 4685 4 vdd
port 46 nsew
rlabel metal3 s 4202 3035 4300 3133 4 vdd
port 46 nsew
rlabel metal3 s 1706 3035 1804 3133 4 vdd
port 46 nsew
rlabel metal3 s 6317 5980 6415 6078 4 vdd
port 46 nsew
rlabel metal3 s 2193 4587 2291 4685 4 vdd
port 46 nsew
rlabel metal3 s 4688 3035 4786 3133 4 vdd
port 46 nsew
rlabel metal3 s 6124 313 6222 411 4 vdd
port 46 nsew
rlabel metal3 s 2766 313 2864 411 4 vdd
port 46 nsew
rlabel metal3 s 5936 3035 6034 3133 4 vdd
port 46 nsew
rlabel metal3 s 1581 4587 1679 4685 4 vdd
port 46 nsew
rlabel metal3 s 1601 5537 1699 5635 4 vdd
port 46 nsew
rlabel metal3 s 1694 2197 1792 2295 4 vdd
port 46 nsew
rlabel metal3 s 4689 4587 4787 4685 4 vdd
port 46 nsew
rlabel metal3 s 3421 5537 3519 5635 4 vdd
port 46 nsew
rlabel metal3 s 4097 5537 4195 5635 4 vdd
port 46 nsew
rlabel metal3 s 4190 2197 4288 2295 4 vdd
port 46 nsew
rlabel metal3 s 2173 5537 2271 5635 4 vdd
port 46 nsew
rlabel metal3 s 5438 2197 5536 2295 4 vdd
port 46 nsew
rlabel metal3 s 6317 7100 6415 7198 4 gnd
port 47 nsew
rlabel metal3 s 5336 4150 5434 4248 4 gnd
port 47 nsew
rlabel metal3 s 5446 4919 5544 5017 4 gnd
port 47 nsew
rlabel metal3 s 2835 5121 2933 5219 4 gnd
port 47 nsew
rlabel metal3 s 4202 3357 4300 3455 4 gnd
port 47 nsew
rlabel metal3 s 1776 1423 1874 1521 4 gnd
port 47 nsew
rlabel metal3 s 4683 5121 4781 5219 4 gnd
port 47 nsew
rlabel metal3 s 4618 1423 4716 1521 4 gnd
port 47 nsew
rlabel metal3 s 1706 3357 1804 3455 4 gnd
port 47 nsew
rlabel metal3 s 5450 3357 5548 3455 4 gnd
port 47 nsew
rlabel metal3 s 2954 3357 3052 3455 4 gnd
port 47 nsew
rlabel metal3 s 5926 4150 6024 4248 4 gnd
port 47 nsew
rlabel metal3 s -49 7100 49 7198 4 gnd
port 47 nsew
rlabel metal3 s 3370 1423 3468 1521 4 gnd
port 47 nsew
rlabel metal3 s 5816 4919 5914 5017 4 gnd
port 47 nsew
rlabel metal3 s 3320 4919 3418 5017 4 gnd
port 47 nsew
rlabel metal3 s 5520 1423 5618 1521 4 gnd
port 47 nsew
rlabel metal3 s 1702 4919 1800 5017 4 gnd
port 47 nsew
rlabel metal3 s 2072 4919 2170 5017 4 gnd
port 47 nsew
rlabel metal3 s 2187 5121 2285 5219 4 gnd
port 47 nsew
rlabel metal3 s 4272 1423 4370 1521 4 gnd
port 47 nsew
rlabel metal3 s 2950 4919 3048 5017 4 gnd
port 47 nsew
rlabel metal3 s 4088 4150 4186 4248 4 gnd
port 47 nsew
rlabel metal3 s 2192 3357 2290 3455 4 gnd
port 47 nsew
rlabel metal3 s 4198 4919 4296 5017 4 gnd
port 47 nsew
rlabel metal3 s 3430 4150 3528 4248 4 gnd
port 47 nsew
rlabel metal3 s 4688 3357 4786 3455 4 gnd
port 47 nsew
rlabel metal3 s 5931 5121 6029 5219 4 gnd
port 47 nsew
rlabel metal3 s 3440 3357 3538 3455 4 gnd
port 47 nsew
rlabel metal3 s 3024 1423 3122 1521 4 gnd
port 47 nsew
rlabel metal3 s 2840 4150 2938 4248 4 gnd
port 47 nsew
rlabel metal3 s 5936 3357 6034 3455 4 gnd
port 47 nsew
rlabel metal3 s 5866 1423 5964 1521 4 gnd
port 47 nsew
rlabel metal3 s 5331 5121 5429 5219 4 gnd
port 47 nsew
rlabel metal3 s 2182 4150 2280 4248 4 gnd
port 47 nsew
rlabel metal3 s 1592 4150 1690 4248 4 gnd
port 47 nsew
rlabel metal3 s 1587 5121 1685 5219 4 gnd
port 47 nsew
rlabel metal3 s 4568 4919 4666 5017 4 gnd
port 47 nsew
rlabel metal3 s 3435 5121 3533 5219 4 gnd
port 47 nsew
rlabel metal3 s 4083 5121 4181 5219 4 gnd
port 47 nsew
rlabel metal3 s 2122 1423 2220 1521 4 gnd
port 47 nsew
rlabel metal3 s 4678 4150 4776 4248 4 gnd
port 47 nsew
<< properties >>
string FIXED_BBOX 0 0 6366 7149
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 795508
string GDS_START 760742
<< end >>
