magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1260 -1260 44720 34384
<< dnwell >>
rect 1758 1760 41740 31384
<< nwell >>
rect 1674 31300 41824 31468
rect 1674 1844 1842 31300
rect 41656 1844 41824 31300
rect 1674 1676 41824 1844
<< nsubdiff >>
rect 2069 31401 2119 31425
rect 2069 31367 2077 31401
rect 2111 31367 2119 31401
rect 2069 31343 2119 31367
rect 2405 31401 2455 31425
rect 2405 31367 2413 31401
rect 2447 31367 2455 31401
rect 2405 31343 2455 31367
rect 2741 31401 2791 31425
rect 2741 31367 2749 31401
rect 2783 31367 2791 31401
rect 2741 31343 2791 31367
rect 3077 31401 3127 31425
rect 3077 31367 3085 31401
rect 3119 31367 3127 31401
rect 3077 31343 3127 31367
rect 3413 31401 3463 31425
rect 3413 31367 3421 31401
rect 3455 31367 3463 31401
rect 3413 31343 3463 31367
rect 3749 31401 3799 31425
rect 3749 31367 3757 31401
rect 3791 31367 3799 31401
rect 3749 31343 3799 31367
rect 4085 31401 4135 31425
rect 4085 31367 4093 31401
rect 4127 31367 4135 31401
rect 4085 31343 4135 31367
rect 4421 31401 4471 31425
rect 4421 31367 4429 31401
rect 4463 31367 4471 31401
rect 4421 31343 4471 31367
rect 4757 31401 4807 31425
rect 4757 31367 4765 31401
rect 4799 31367 4807 31401
rect 4757 31343 4807 31367
rect 5093 31401 5143 31425
rect 5093 31367 5101 31401
rect 5135 31367 5143 31401
rect 5093 31343 5143 31367
rect 5429 31401 5479 31425
rect 5429 31367 5437 31401
rect 5471 31367 5479 31401
rect 5429 31343 5479 31367
rect 5765 31401 5815 31425
rect 5765 31367 5773 31401
rect 5807 31367 5815 31401
rect 5765 31343 5815 31367
rect 6101 31401 6151 31425
rect 6101 31367 6109 31401
rect 6143 31367 6151 31401
rect 6101 31343 6151 31367
rect 6437 31401 6487 31425
rect 6437 31367 6445 31401
rect 6479 31367 6487 31401
rect 6437 31343 6487 31367
rect 6773 31401 6823 31425
rect 6773 31367 6781 31401
rect 6815 31367 6823 31401
rect 6773 31343 6823 31367
rect 7109 31401 7159 31425
rect 7109 31367 7117 31401
rect 7151 31367 7159 31401
rect 7109 31343 7159 31367
rect 7445 31401 7495 31425
rect 7445 31367 7453 31401
rect 7487 31367 7495 31401
rect 7445 31343 7495 31367
rect 7781 31401 7831 31425
rect 7781 31367 7789 31401
rect 7823 31367 7831 31401
rect 7781 31343 7831 31367
rect 8117 31401 8167 31425
rect 8117 31367 8125 31401
rect 8159 31367 8167 31401
rect 8117 31343 8167 31367
rect 8453 31401 8503 31425
rect 8453 31367 8461 31401
rect 8495 31367 8503 31401
rect 8453 31343 8503 31367
rect 8789 31401 8839 31425
rect 8789 31367 8797 31401
rect 8831 31367 8839 31401
rect 8789 31343 8839 31367
rect 9125 31401 9175 31425
rect 9125 31367 9133 31401
rect 9167 31367 9175 31401
rect 9125 31343 9175 31367
rect 9461 31401 9511 31425
rect 9461 31367 9469 31401
rect 9503 31367 9511 31401
rect 9461 31343 9511 31367
rect 9797 31401 9847 31425
rect 9797 31367 9805 31401
rect 9839 31367 9847 31401
rect 9797 31343 9847 31367
rect 10133 31401 10183 31425
rect 10133 31367 10141 31401
rect 10175 31367 10183 31401
rect 10133 31343 10183 31367
rect 10469 31401 10519 31425
rect 10469 31367 10477 31401
rect 10511 31367 10519 31401
rect 10469 31343 10519 31367
rect 10805 31401 10855 31425
rect 10805 31367 10813 31401
rect 10847 31367 10855 31401
rect 10805 31343 10855 31367
rect 11141 31401 11191 31425
rect 11141 31367 11149 31401
rect 11183 31367 11191 31401
rect 11141 31343 11191 31367
rect 11477 31401 11527 31425
rect 11477 31367 11485 31401
rect 11519 31367 11527 31401
rect 11477 31343 11527 31367
rect 11813 31401 11863 31425
rect 11813 31367 11821 31401
rect 11855 31367 11863 31401
rect 11813 31343 11863 31367
rect 12149 31401 12199 31425
rect 12149 31367 12157 31401
rect 12191 31367 12199 31401
rect 12149 31343 12199 31367
rect 12485 31401 12535 31425
rect 12485 31367 12493 31401
rect 12527 31367 12535 31401
rect 12485 31343 12535 31367
rect 12821 31401 12871 31425
rect 12821 31367 12829 31401
rect 12863 31367 12871 31401
rect 12821 31343 12871 31367
rect 13157 31401 13207 31425
rect 13157 31367 13165 31401
rect 13199 31367 13207 31401
rect 13157 31343 13207 31367
rect 13493 31401 13543 31425
rect 13493 31367 13501 31401
rect 13535 31367 13543 31401
rect 13493 31343 13543 31367
rect 13829 31401 13879 31425
rect 13829 31367 13837 31401
rect 13871 31367 13879 31401
rect 13829 31343 13879 31367
rect 14165 31401 14215 31425
rect 14165 31367 14173 31401
rect 14207 31367 14215 31401
rect 14165 31343 14215 31367
rect 14501 31401 14551 31425
rect 14501 31367 14509 31401
rect 14543 31367 14551 31401
rect 14501 31343 14551 31367
rect 14837 31401 14887 31425
rect 14837 31367 14845 31401
rect 14879 31367 14887 31401
rect 14837 31343 14887 31367
rect 15173 31401 15223 31425
rect 15173 31367 15181 31401
rect 15215 31367 15223 31401
rect 15173 31343 15223 31367
rect 15509 31401 15559 31425
rect 15509 31367 15517 31401
rect 15551 31367 15559 31401
rect 15509 31343 15559 31367
rect 15845 31401 15895 31425
rect 15845 31367 15853 31401
rect 15887 31367 15895 31401
rect 15845 31343 15895 31367
rect 16181 31401 16231 31425
rect 16181 31367 16189 31401
rect 16223 31367 16231 31401
rect 16181 31343 16231 31367
rect 16517 31401 16567 31425
rect 16517 31367 16525 31401
rect 16559 31367 16567 31401
rect 16517 31343 16567 31367
rect 16853 31401 16903 31425
rect 16853 31367 16861 31401
rect 16895 31367 16903 31401
rect 16853 31343 16903 31367
rect 17189 31401 17239 31425
rect 17189 31367 17197 31401
rect 17231 31367 17239 31401
rect 17189 31343 17239 31367
rect 17525 31401 17575 31425
rect 17525 31367 17533 31401
rect 17567 31367 17575 31401
rect 17525 31343 17575 31367
rect 17861 31401 17911 31425
rect 17861 31367 17869 31401
rect 17903 31367 17911 31401
rect 17861 31343 17911 31367
rect 18197 31401 18247 31425
rect 18197 31367 18205 31401
rect 18239 31367 18247 31401
rect 18197 31343 18247 31367
rect 18533 31401 18583 31425
rect 18533 31367 18541 31401
rect 18575 31367 18583 31401
rect 18533 31343 18583 31367
rect 18869 31401 18919 31425
rect 18869 31367 18877 31401
rect 18911 31367 18919 31401
rect 18869 31343 18919 31367
rect 19205 31401 19255 31425
rect 19205 31367 19213 31401
rect 19247 31367 19255 31401
rect 19205 31343 19255 31367
rect 19541 31401 19591 31425
rect 19541 31367 19549 31401
rect 19583 31367 19591 31401
rect 19541 31343 19591 31367
rect 19877 31401 19927 31425
rect 19877 31367 19885 31401
rect 19919 31367 19927 31401
rect 19877 31343 19927 31367
rect 20213 31401 20263 31425
rect 20213 31367 20221 31401
rect 20255 31367 20263 31401
rect 20213 31343 20263 31367
rect 20549 31401 20599 31425
rect 20549 31367 20557 31401
rect 20591 31367 20599 31401
rect 20549 31343 20599 31367
rect 20885 31401 20935 31425
rect 20885 31367 20893 31401
rect 20927 31367 20935 31401
rect 20885 31343 20935 31367
rect 21221 31401 21271 31425
rect 21221 31367 21229 31401
rect 21263 31367 21271 31401
rect 21221 31343 21271 31367
rect 21557 31401 21607 31425
rect 21557 31367 21565 31401
rect 21599 31367 21607 31401
rect 21557 31343 21607 31367
rect 21893 31401 21943 31425
rect 21893 31367 21901 31401
rect 21935 31367 21943 31401
rect 21893 31343 21943 31367
rect 22229 31401 22279 31425
rect 22229 31367 22237 31401
rect 22271 31367 22279 31401
rect 22229 31343 22279 31367
rect 22565 31401 22615 31425
rect 22565 31367 22573 31401
rect 22607 31367 22615 31401
rect 22565 31343 22615 31367
rect 22901 31401 22951 31425
rect 22901 31367 22909 31401
rect 22943 31367 22951 31401
rect 22901 31343 22951 31367
rect 23237 31401 23287 31425
rect 23237 31367 23245 31401
rect 23279 31367 23287 31401
rect 23237 31343 23287 31367
rect 23573 31401 23623 31425
rect 23573 31367 23581 31401
rect 23615 31367 23623 31401
rect 23573 31343 23623 31367
rect 23909 31401 23959 31425
rect 23909 31367 23917 31401
rect 23951 31367 23959 31401
rect 23909 31343 23959 31367
rect 24245 31401 24295 31425
rect 24245 31367 24253 31401
rect 24287 31367 24295 31401
rect 24245 31343 24295 31367
rect 24581 31401 24631 31425
rect 24581 31367 24589 31401
rect 24623 31367 24631 31401
rect 24581 31343 24631 31367
rect 24917 31401 24967 31425
rect 24917 31367 24925 31401
rect 24959 31367 24967 31401
rect 24917 31343 24967 31367
rect 25253 31401 25303 31425
rect 25253 31367 25261 31401
rect 25295 31367 25303 31401
rect 25253 31343 25303 31367
rect 25589 31401 25639 31425
rect 25589 31367 25597 31401
rect 25631 31367 25639 31401
rect 25589 31343 25639 31367
rect 25925 31401 25975 31425
rect 25925 31367 25933 31401
rect 25967 31367 25975 31401
rect 25925 31343 25975 31367
rect 26261 31401 26311 31425
rect 26261 31367 26269 31401
rect 26303 31367 26311 31401
rect 26261 31343 26311 31367
rect 26597 31401 26647 31425
rect 26597 31367 26605 31401
rect 26639 31367 26647 31401
rect 26597 31343 26647 31367
rect 26933 31401 26983 31425
rect 26933 31367 26941 31401
rect 26975 31367 26983 31401
rect 26933 31343 26983 31367
rect 27269 31401 27319 31425
rect 27269 31367 27277 31401
rect 27311 31367 27319 31401
rect 27269 31343 27319 31367
rect 27605 31401 27655 31425
rect 27605 31367 27613 31401
rect 27647 31367 27655 31401
rect 27605 31343 27655 31367
rect 27941 31401 27991 31425
rect 27941 31367 27949 31401
rect 27983 31367 27991 31401
rect 27941 31343 27991 31367
rect 28277 31401 28327 31425
rect 28277 31367 28285 31401
rect 28319 31367 28327 31401
rect 28277 31343 28327 31367
rect 28613 31401 28663 31425
rect 28613 31367 28621 31401
rect 28655 31367 28663 31401
rect 28613 31343 28663 31367
rect 28949 31401 28999 31425
rect 28949 31367 28957 31401
rect 28991 31367 28999 31401
rect 28949 31343 28999 31367
rect 29285 31401 29335 31425
rect 29285 31367 29293 31401
rect 29327 31367 29335 31401
rect 29285 31343 29335 31367
rect 29621 31401 29671 31425
rect 29621 31367 29629 31401
rect 29663 31367 29671 31401
rect 29621 31343 29671 31367
rect 29957 31401 30007 31425
rect 29957 31367 29965 31401
rect 29999 31367 30007 31401
rect 29957 31343 30007 31367
rect 30293 31401 30343 31425
rect 30293 31367 30301 31401
rect 30335 31367 30343 31401
rect 30293 31343 30343 31367
rect 30629 31401 30679 31425
rect 30629 31367 30637 31401
rect 30671 31367 30679 31401
rect 30629 31343 30679 31367
rect 30965 31401 31015 31425
rect 30965 31367 30973 31401
rect 31007 31367 31015 31401
rect 30965 31343 31015 31367
rect 31301 31401 31351 31425
rect 31301 31367 31309 31401
rect 31343 31367 31351 31401
rect 31301 31343 31351 31367
rect 31637 31401 31687 31425
rect 31637 31367 31645 31401
rect 31679 31367 31687 31401
rect 31637 31343 31687 31367
rect 31973 31401 32023 31425
rect 31973 31367 31981 31401
rect 32015 31367 32023 31401
rect 31973 31343 32023 31367
rect 32309 31401 32359 31425
rect 32309 31367 32317 31401
rect 32351 31367 32359 31401
rect 32309 31343 32359 31367
rect 32645 31401 32695 31425
rect 32645 31367 32653 31401
rect 32687 31367 32695 31401
rect 32645 31343 32695 31367
rect 32981 31401 33031 31425
rect 32981 31367 32989 31401
rect 33023 31367 33031 31401
rect 32981 31343 33031 31367
rect 33317 31401 33367 31425
rect 33317 31367 33325 31401
rect 33359 31367 33367 31401
rect 33317 31343 33367 31367
rect 33653 31401 33703 31425
rect 33653 31367 33661 31401
rect 33695 31367 33703 31401
rect 33653 31343 33703 31367
rect 33989 31401 34039 31425
rect 33989 31367 33997 31401
rect 34031 31367 34039 31401
rect 33989 31343 34039 31367
rect 34325 31401 34375 31425
rect 34325 31367 34333 31401
rect 34367 31367 34375 31401
rect 34325 31343 34375 31367
rect 34661 31401 34711 31425
rect 34661 31367 34669 31401
rect 34703 31367 34711 31401
rect 34661 31343 34711 31367
rect 34997 31401 35047 31425
rect 34997 31367 35005 31401
rect 35039 31367 35047 31401
rect 34997 31343 35047 31367
rect 35333 31401 35383 31425
rect 35333 31367 35341 31401
rect 35375 31367 35383 31401
rect 35333 31343 35383 31367
rect 35669 31401 35719 31425
rect 35669 31367 35677 31401
rect 35711 31367 35719 31401
rect 35669 31343 35719 31367
rect 36005 31401 36055 31425
rect 36005 31367 36013 31401
rect 36047 31367 36055 31401
rect 36005 31343 36055 31367
rect 36341 31401 36391 31425
rect 36341 31367 36349 31401
rect 36383 31367 36391 31401
rect 36341 31343 36391 31367
rect 36677 31401 36727 31425
rect 36677 31367 36685 31401
rect 36719 31367 36727 31401
rect 36677 31343 36727 31367
rect 37013 31401 37063 31425
rect 37013 31367 37021 31401
rect 37055 31367 37063 31401
rect 37013 31343 37063 31367
rect 37349 31401 37399 31425
rect 37349 31367 37357 31401
rect 37391 31367 37399 31401
rect 37349 31343 37399 31367
rect 37685 31401 37735 31425
rect 37685 31367 37693 31401
rect 37727 31367 37735 31401
rect 37685 31343 37735 31367
rect 38021 31401 38071 31425
rect 38021 31367 38029 31401
rect 38063 31367 38071 31401
rect 38021 31343 38071 31367
rect 38357 31401 38407 31425
rect 38357 31367 38365 31401
rect 38399 31367 38407 31401
rect 38357 31343 38407 31367
rect 38693 31401 38743 31425
rect 38693 31367 38701 31401
rect 38735 31367 38743 31401
rect 38693 31343 38743 31367
rect 39029 31401 39079 31425
rect 39029 31367 39037 31401
rect 39071 31367 39079 31401
rect 39029 31343 39079 31367
rect 39365 31401 39415 31425
rect 39365 31367 39373 31401
rect 39407 31367 39415 31401
rect 39365 31343 39415 31367
rect 39701 31401 39751 31425
rect 39701 31367 39709 31401
rect 39743 31367 39751 31401
rect 39701 31343 39751 31367
rect 40037 31401 40087 31425
rect 40037 31367 40045 31401
rect 40079 31367 40087 31401
rect 40037 31343 40087 31367
rect 40373 31401 40423 31425
rect 40373 31367 40381 31401
rect 40415 31367 40423 31401
rect 40373 31343 40423 31367
rect 40709 31401 40759 31425
rect 40709 31367 40717 31401
rect 40751 31367 40759 31401
rect 40709 31343 40759 31367
rect 41045 31401 41095 31425
rect 41045 31367 41053 31401
rect 41087 31367 41095 31401
rect 41045 31343 41095 31367
rect 1733 31009 1783 31033
rect 1733 30975 1741 31009
rect 1775 30975 1783 31009
rect 1733 30951 1783 30975
rect 41715 31009 41765 31033
rect 41715 30975 41723 31009
rect 41757 30975 41765 31009
rect 41715 30951 41765 30975
rect 1733 30673 1783 30697
rect 1733 30639 1741 30673
rect 1775 30639 1783 30673
rect 1733 30615 1783 30639
rect 41715 30673 41765 30697
rect 41715 30639 41723 30673
rect 41757 30639 41765 30673
rect 41715 30615 41765 30639
rect 1733 30337 1783 30361
rect 1733 30303 1741 30337
rect 1775 30303 1783 30337
rect 1733 30279 1783 30303
rect 41715 30337 41765 30361
rect 41715 30303 41723 30337
rect 41757 30303 41765 30337
rect 41715 30279 41765 30303
rect 1733 30001 1783 30025
rect 1733 29967 1741 30001
rect 1775 29967 1783 30001
rect 1733 29943 1783 29967
rect 41715 30001 41765 30025
rect 41715 29967 41723 30001
rect 41757 29967 41765 30001
rect 41715 29943 41765 29967
rect 1733 29665 1783 29689
rect 1733 29631 1741 29665
rect 1775 29631 1783 29665
rect 1733 29607 1783 29631
rect 41715 29665 41765 29689
rect 41715 29631 41723 29665
rect 41757 29631 41765 29665
rect 41715 29607 41765 29631
rect 1733 29329 1783 29353
rect 1733 29295 1741 29329
rect 1775 29295 1783 29329
rect 1733 29271 1783 29295
rect 41715 29329 41765 29353
rect 41715 29295 41723 29329
rect 41757 29295 41765 29329
rect 41715 29271 41765 29295
rect 1733 28993 1783 29017
rect 1733 28959 1741 28993
rect 1775 28959 1783 28993
rect 1733 28935 1783 28959
rect 41715 28993 41765 29017
rect 41715 28959 41723 28993
rect 41757 28959 41765 28993
rect 41715 28935 41765 28959
rect 1733 28657 1783 28681
rect 1733 28623 1741 28657
rect 1775 28623 1783 28657
rect 1733 28599 1783 28623
rect 41715 28657 41765 28681
rect 41715 28623 41723 28657
rect 41757 28623 41765 28657
rect 41715 28599 41765 28623
rect 1733 28321 1783 28345
rect 1733 28287 1741 28321
rect 1775 28287 1783 28321
rect 1733 28263 1783 28287
rect 41715 28321 41765 28345
rect 41715 28287 41723 28321
rect 41757 28287 41765 28321
rect 41715 28263 41765 28287
rect 1733 27985 1783 28009
rect 1733 27951 1741 27985
rect 1775 27951 1783 27985
rect 1733 27927 1783 27951
rect 41715 27985 41765 28009
rect 41715 27951 41723 27985
rect 41757 27951 41765 27985
rect 41715 27927 41765 27951
rect 1733 27649 1783 27673
rect 1733 27615 1741 27649
rect 1775 27615 1783 27649
rect 1733 27591 1783 27615
rect 41715 27649 41765 27673
rect 41715 27615 41723 27649
rect 41757 27615 41765 27649
rect 41715 27591 41765 27615
rect 1733 27313 1783 27337
rect 1733 27279 1741 27313
rect 1775 27279 1783 27313
rect 1733 27255 1783 27279
rect 41715 27313 41765 27337
rect 41715 27279 41723 27313
rect 41757 27279 41765 27313
rect 41715 27255 41765 27279
rect 1733 26977 1783 27001
rect 1733 26943 1741 26977
rect 1775 26943 1783 26977
rect 1733 26919 1783 26943
rect 41715 26977 41765 27001
rect 41715 26943 41723 26977
rect 41757 26943 41765 26977
rect 41715 26919 41765 26943
rect 1733 26641 1783 26665
rect 1733 26607 1741 26641
rect 1775 26607 1783 26641
rect 1733 26583 1783 26607
rect 41715 26641 41765 26665
rect 41715 26607 41723 26641
rect 41757 26607 41765 26641
rect 41715 26583 41765 26607
rect 1733 26305 1783 26329
rect 1733 26271 1741 26305
rect 1775 26271 1783 26305
rect 1733 26247 1783 26271
rect 41715 26305 41765 26329
rect 41715 26271 41723 26305
rect 41757 26271 41765 26305
rect 41715 26247 41765 26271
rect 1733 25969 1783 25993
rect 1733 25935 1741 25969
rect 1775 25935 1783 25969
rect 1733 25911 1783 25935
rect 41715 25969 41765 25993
rect 41715 25935 41723 25969
rect 41757 25935 41765 25969
rect 41715 25911 41765 25935
rect 1733 25633 1783 25657
rect 1733 25599 1741 25633
rect 1775 25599 1783 25633
rect 1733 25575 1783 25599
rect 41715 25633 41765 25657
rect 41715 25599 41723 25633
rect 41757 25599 41765 25633
rect 41715 25575 41765 25599
rect 1733 25297 1783 25321
rect 1733 25263 1741 25297
rect 1775 25263 1783 25297
rect 1733 25239 1783 25263
rect 41715 25297 41765 25321
rect 41715 25263 41723 25297
rect 41757 25263 41765 25297
rect 41715 25239 41765 25263
rect 1733 24961 1783 24985
rect 1733 24927 1741 24961
rect 1775 24927 1783 24961
rect 1733 24903 1783 24927
rect 41715 24961 41765 24985
rect 41715 24927 41723 24961
rect 41757 24927 41765 24961
rect 41715 24903 41765 24927
rect 1733 24625 1783 24649
rect 1733 24591 1741 24625
rect 1775 24591 1783 24625
rect 1733 24567 1783 24591
rect 41715 24625 41765 24649
rect 41715 24591 41723 24625
rect 41757 24591 41765 24625
rect 41715 24567 41765 24591
rect 1733 24289 1783 24313
rect 1733 24255 1741 24289
rect 1775 24255 1783 24289
rect 1733 24231 1783 24255
rect 41715 24289 41765 24313
rect 41715 24255 41723 24289
rect 41757 24255 41765 24289
rect 41715 24231 41765 24255
rect 1733 23953 1783 23977
rect 1733 23919 1741 23953
rect 1775 23919 1783 23953
rect 1733 23895 1783 23919
rect 41715 23953 41765 23977
rect 41715 23919 41723 23953
rect 41757 23919 41765 23953
rect 41715 23895 41765 23919
rect 1733 23617 1783 23641
rect 1733 23583 1741 23617
rect 1775 23583 1783 23617
rect 1733 23559 1783 23583
rect 41715 23617 41765 23641
rect 41715 23583 41723 23617
rect 41757 23583 41765 23617
rect 41715 23559 41765 23583
rect 1733 23281 1783 23305
rect 1733 23247 1741 23281
rect 1775 23247 1783 23281
rect 1733 23223 1783 23247
rect 41715 23281 41765 23305
rect 41715 23247 41723 23281
rect 41757 23247 41765 23281
rect 41715 23223 41765 23247
rect 1733 22945 1783 22969
rect 1733 22911 1741 22945
rect 1775 22911 1783 22945
rect 1733 22887 1783 22911
rect 41715 22945 41765 22969
rect 41715 22911 41723 22945
rect 41757 22911 41765 22945
rect 41715 22887 41765 22911
rect 1733 22609 1783 22633
rect 1733 22575 1741 22609
rect 1775 22575 1783 22609
rect 1733 22551 1783 22575
rect 41715 22609 41765 22633
rect 41715 22575 41723 22609
rect 41757 22575 41765 22609
rect 41715 22551 41765 22575
rect 1733 22273 1783 22297
rect 1733 22239 1741 22273
rect 1775 22239 1783 22273
rect 1733 22215 1783 22239
rect 41715 22273 41765 22297
rect 41715 22239 41723 22273
rect 41757 22239 41765 22273
rect 41715 22215 41765 22239
rect 1733 21937 1783 21961
rect 1733 21903 1741 21937
rect 1775 21903 1783 21937
rect 1733 21879 1783 21903
rect 41715 21937 41765 21961
rect 41715 21903 41723 21937
rect 41757 21903 41765 21937
rect 41715 21879 41765 21903
rect 1733 21601 1783 21625
rect 1733 21567 1741 21601
rect 1775 21567 1783 21601
rect 1733 21543 1783 21567
rect 41715 21601 41765 21625
rect 41715 21567 41723 21601
rect 41757 21567 41765 21601
rect 41715 21543 41765 21567
rect 1733 21265 1783 21289
rect 1733 21231 1741 21265
rect 1775 21231 1783 21265
rect 1733 21207 1783 21231
rect 41715 21265 41765 21289
rect 41715 21231 41723 21265
rect 41757 21231 41765 21265
rect 41715 21207 41765 21231
rect 1733 20929 1783 20953
rect 1733 20895 1741 20929
rect 1775 20895 1783 20929
rect 1733 20871 1783 20895
rect 41715 20929 41765 20953
rect 41715 20895 41723 20929
rect 41757 20895 41765 20929
rect 41715 20871 41765 20895
rect 1733 20593 1783 20617
rect 1733 20559 1741 20593
rect 1775 20559 1783 20593
rect 1733 20535 1783 20559
rect 41715 20593 41765 20617
rect 41715 20559 41723 20593
rect 41757 20559 41765 20593
rect 41715 20535 41765 20559
rect 1733 20257 1783 20281
rect 1733 20223 1741 20257
rect 1775 20223 1783 20257
rect 1733 20199 1783 20223
rect 41715 20257 41765 20281
rect 41715 20223 41723 20257
rect 41757 20223 41765 20257
rect 41715 20199 41765 20223
rect 1733 19921 1783 19945
rect 1733 19887 1741 19921
rect 1775 19887 1783 19921
rect 1733 19863 1783 19887
rect 41715 19921 41765 19945
rect 41715 19887 41723 19921
rect 41757 19887 41765 19921
rect 41715 19863 41765 19887
rect 1733 19585 1783 19609
rect 1733 19551 1741 19585
rect 1775 19551 1783 19585
rect 1733 19527 1783 19551
rect 41715 19585 41765 19609
rect 41715 19551 41723 19585
rect 41757 19551 41765 19585
rect 41715 19527 41765 19551
rect 1733 19249 1783 19273
rect 1733 19215 1741 19249
rect 1775 19215 1783 19249
rect 1733 19191 1783 19215
rect 41715 19249 41765 19273
rect 41715 19215 41723 19249
rect 41757 19215 41765 19249
rect 41715 19191 41765 19215
rect 1733 18913 1783 18937
rect 1733 18879 1741 18913
rect 1775 18879 1783 18913
rect 1733 18855 1783 18879
rect 41715 18913 41765 18937
rect 41715 18879 41723 18913
rect 41757 18879 41765 18913
rect 41715 18855 41765 18879
rect 1733 18577 1783 18601
rect 1733 18543 1741 18577
rect 1775 18543 1783 18577
rect 1733 18519 1783 18543
rect 41715 18577 41765 18601
rect 41715 18543 41723 18577
rect 41757 18543 41765 18577
rect 41715 18519 41765 18543
rect 1733 18241 1783 18265
rect 1733 18207 1741 18241
rect 1775 18207 1783 18241
rect 1733 18183 1783 18207
rect 41715 18241 41765 18265
rect 41715 18207 41723 18241
rect 41757 18207 41765 18241
rect 41715 18183 41765 18207
rect 1733 17905 1783 17929
rect 1733 17871 1741 17905
rect 1775 17871 1783 17905
rect 1733 17847 1783 17871
rect 41715 17905 41765 17929
rect 41715 17871 41723 17905
rect 41757 17871 41765 17905
rect 41715 17847 41765 17871
rect 1733 17569 1783 17593
rect 1733 17535 1741 17569
rect 1775 17535 1783 17569
rect 1733 17511 1783 17535
rect 41715 17569 41765 17593
rect 41715 17535 41723 17569
rect 41757 17535 41765 17569
rect 41715 17511 41765 17535
rect 1733 17233 1783 17257
rect 1733 17199 1741 17233
rect 1775 17199 1783 17233
rect 1733 17175 1783 17199
rect 41715 17233 41765 17257
rect 41715 17199 41723 17233
rect 41757 17199 41765 17233
rect 41715 17175 41765 17199
rect 1733 16897 1783 16921
rect 1733 16863 1741 16897
rect 1775 16863 1783 16897
rect 1733 16839 1783 16863
rect 41715 16897 41765 16921
rect 41715 16863 41723 16897
rect 41757 16863 41765 16897
rect 41715 16839 41765 16863
rect 1733 16561 1783 16585
rect 1733 16527 1741 16561
rect 1775 16527 1783 16561
rect 1733 16503 1783 16527
rect 41715 16561 41765 16585
rect 41715 16527 41723 16561
rect 41757 16527 41765 16561
rect 41715 16503 41765 16527
rect 1733 16225 1783 16249
rect 1733 16191 1741 16225
rect 1775 16191 1783 16225
rect 1733 16167 1783 16191
rect 41715 16225 41765 16249
rect 41715 16191 41723 16225
rect 41757 16191 41765 16225
rect 41715 16167 41765 16191
rect 1733 15889 1783 15913
rect 1733 15855 1741 15889
rect 1775 15855 1783 15889
rect 1733 15831 1783 15855
rect 41715 15889 41765 15913
rect 41715 15855 41723 15889
rect 41757 15855 41765 15889
rect 41715 15831 41765 15855
rect 1733 15553 1783 15577
rect 1733 15519 1741 15553
rect 1775 15519 1783 15553
rect 1733 15495 1783 15519
rect 41715 15553 41765 15577
rect 41715 15519 41723 15553
rect 41757 15519 41765 15553
rect 41715 15495 41765 15519
rect 1733 15217 1783 15241
rect 1733 15183 1741 15217
rect 1775 15183 1783 15217
rect 1733 15159 1783 15183
rect 41715 15217 41765 15241
rect 41715 15183 41723 15217
rect 41757 15183 41765 15217
rect 41715 15159 41765 15183
rect 1733 14881 1783 14905
rect 1733 14847 1741 14881
rect 1775 14847 1783 14881
rect 1733 14823 1783 14847
rect 41715 14881 41765 14905
rect 41715 14847 41723 14881
rect 41757 14847 41765 14881
rect 41715 14823 41765 14847
rect 1733 14545 1783 14569
rect 1733 14511 1741 14545
rect 1775 14511 1783 14545
rect 1733 14487 1783 14511
rect 41715 14545 41765 14569
rect 41715 14511 41723 14545
rect 41757 14511 41765 14545
rect 41715 14487 41765 14511
rect 1733 14209 1783 14233
rect 1733 14175 1741 14209
rect 1775 14175 1783 14209
rect 1733 14151 1783 14175
rect 41715 14209 41765 14233
rect 41715 14175 41723 14209
rect 41757 14175 41765 14209
rect 41715 14151 41765 14175
rect 1733 13873 1783 13897
rect 1733 13839 1741 13873
rect 1775 13839 1783 13873
rect 1733 13815 1783 13839
rect 41715 13873 41765 13897
rect 41715 13839 41723 13873
rect 41757 13839 41765 13873
rect 41715 13815 41765 13839
rect 1733 13537 1783 13561
rect 1733 13503 1741 13537
rect 1775 13503 1783 13537
rect 1733 13479 1783 13503
rect 41715 13537 41765 13561
rect 41715 13503 41723 13537
rect 41757 13503 41765 13537
rect 41715 13479 41765 13503
rect 1733 13201 1783 13225
rect 1733 13167 1741 13201
rect 1775 13167 1783 13201
rect 1733 13143 1783 13167
rect 41715 13201 41765 13225
rect 41715 13167 41723 13201
rect 41757 13167 41765 13201
rect 41715 13143 41765 13167
rect 1733 12865 1783 12889
rect 1733 12831 1741 12865
rect 1775 12831 1783 12865
rect 1733 12807 1783 12831
rect 41715 12865 41765 12889
rect 41715 12831 41723 12865
rect 41757 12831 41765 12865
rect 41715 12807 41765 12831
rect 1733 12529 1783 12553
rect 1733 12495 1741 12529
rect 1775 12495 1783 12529
rect 1733 12471 1783 12495
rect 41715 12529 41765 12553
rect 41715 12495 41723 12529
rect 41757 12495 41765 12529
rect 41715 12471 41765 12495
rect 1733 12193 1783 12217
rect 1733 12159 1741 12193
rect 1775 12159 1783 12193
rect 1733 12135 1783 12159
rect 41715 12193 41765 12217
rect 41715 12159 41723 12193
rect 41757 12159 41765 12193
rect 41715 12135 41765 12159
rect 1733 11857 1783 11881
rect 1733 11823 1741 11857
rect 1775 11823 1783 11857
rect 1733 11799 1783 11823
rect 41715 11857 41765 11881
rect 41715 11823 41723 11857
rect 41757 11823 41765 11857
rect 41715 11799 41765 11823
rect 1733 11521 1783 11545
rect 1733 11487 1741 11521
rect 1775 11487 1783 11521
rect 1733 11463 1783 11487
rect 41715 11521 41765 11545
rect 41715 11487 41723 11521
rect 41757 11487 41765 11521
rect 41715 11463 41765 11487
rect 1733 11185 1783 11209
rect 1733 11151 1741 11185
rect 1775 11151 1783 11185
rect 1733 11127 1783 11151
rect 41715 11185 41765 11209
rect 41715 11151 41723 11185
rect 41757 11151 41765 11185
rect 41715 11127 41765 11151
rect 1733 10849 1783 10873
rect 1733 10815 1741 10849
rect 1775 10815 1783 10849
rect 1733 10791 1783 10815
rect 41715 10849 41765 10873
rect 41715 10815 41723 10849
rect 41757 10815 41765 10849
rect 41715 10791 41765 10815
rect 1733 10513 1783 10537
rect 1733 10479 1741 10513
rect 1775 10479 1783 10513
rect 1733 10455 1783 10479
rect 41715 10513 41765 10537
rect 41715 10479 41723 10513
rect 41757 10479 41765 10513
rect 41715 10455 41765 10479
rect 1733 10177 1783 10201
rect 1733 10143 1741 10177
rect 1775 10143 1783 10177
rect 1733 10119 1783 10143
rect 41715 10177 41765 10201
rect 41715 10143 41723 10177
rect 41757 10143 41765 10177
rect 41715 10119 41765 10143
rect 1733 9841 1783 9865
rect 1733 9807 1741 9841
rect 1775 9807 1783 9841
rect 1733 9783 1783 9807
rect 41715 9841 41765 9865
rect 41715 9807 41723 9841
rect 41757 9807 41765 9841
rect 41715 9783 41765 9807
rect 1733 9505 1783 9529
rect 1733 9471 1741 9505
rect 1775 9471 1783 9505
rect 1733 9447 1783 9471
rect 41715 9505 41765 9529
rect 41715 9471 41723 9505
rect 41757 9471 41765 9505
rect 41715 9447 41765 9471
rect 1733 9169 1783 9193
rect 1733 9135 1741 9169
rect 1775 9135 1783 9169
rect 1733 9111 1783 9135
rect 41715 9169 41765 9193
rect 41715 9135 41723 9169
rect 41757 9135 41765 9169
rect 41715 9111 41765 9135
rect 1733 8833 1783 8857
rect 1733 8799 1741 8833
rect 1775 8799 1783 8833
rect 1733 8775 1783 8799
rect 41715 8833 41765 8857
rect 41715 8799 41723 8833
rect 41757 8799 41765 8833
rect 41715 8775 41765 8799
rect 1733 8497 1783 8521
rect 1733 8463 1741 8497
rect 1775 8463 1783 8497
rect 1733 8439 1783 8463
rect 41715 8497 41765 8521
rect 41715 8463 41723 8497
rect 41757 8463 41765 8497
rect 41715 8439 41765 8463
rect 1733 8161 1783 8185
rect 1733 8127 1741 8161
rect 1775 8127 1783 8161
rect 1733 8103 1783 8127
rect 41715 8161 41765 8185
rect 41715 8127 41723 8161
rect 41757 8127 41765 8161
rect 41715 8103 41765 8127
rect 1733 7825 1783 7849
rect 1733 7791 1741 7825
rect 1775 7791 1783 7825
rect 1733 7767 1783 7791
rect 41715 7825 41765 7849
rect 41715 7791 41723 7825
rect 41757 7791 41765 7825
rect 41715 7767 41765 7791
rect 1733 7489 1783 7513
rect 1733 7455 1741 7489
rect 1775 7455 1783 7489
rect 1733 7431 1783 7455
rect 41715 7489 41765 7513
rect 41715 7455 41723 7489
rect 41757 7455 41765 7489
rect 41715 7431 41765 7455
rect 1733 7153 1783 7177
rect 1733 7119 1741 7153
rect 1775 7119 1783 7153
rect 1733 7095 1783 7119
rect 41715 7153 41765 7177
rect 41715 7119 41723 7153
rect 41757 7119 41765 7153
rect 41715 7095 41765 7119
rect 1733 6817 1783 6841
rect 1733 6783 1741 6817
rect 1775 6783 1783 6817
rect 1733 6759 1783 6783
rect 41715 6817 41765 6841
rect 41715 6783 41723 6817
rect 41757 6783 41765 6817
rect 41715 6759 41765 6783
rect 1733 6481 1783 6505
rect 1733 6447 1741 6481
rect 1775 6447 1783 6481
rect 1733 6423 1783 6447
rect 41715 6481 41765 6505
rect 41715 6447 41723 6481
rect 41757 6447 41765 6481
rect 41715 6423 41765 6447
rect 1733 6145 1783 6169
rect 1733 6111 1741 6145
rect 1775 6111 1783 6145
rect 1733 6087 1783 6111
rect 41715 6145 41765 6169
rect 41715 6111 41723 6145
rect 41757 6111 41765 6145
rect 41715 6087 41765 6111
rect 1733 5809 1783 5833
rect 1733 5775 1741 5809
rect 1775 5775 1783 5809
rect 1733 5751 1783 5775
rect 41715 5809 41765 5833
rect 41715 5775 41723 5809
rect 41757 5775 41765 5809
rect 41715 5751 41765 5775
rect 1733 5473 1783 5497
rect 1733 5439 1741 5473
rect 1775 5439 1783 5473
rect 1733 5415 1783 5439
rect 41715 5473 41765 5497
rect 41715 5439 41723 5473
rect 41757 5439 41765 5473
rect 41715 5415 41765 5439
rect 1733 5137 1783 5161
rect 1733 5103 1741 5137
rect 1775 5103 1783 5137
rect 1733 5079 1783 5103
rect 41715 5137 41765 5161
rect 41715 5103 41723 5137
rect 41757 5103 41765 5137
rect 41715 5079 41765 5103
rect 1733 4801 1783 4825
rect 1733 4767 1741 4801
rect 1775 4767 1783 4801
rect 1733 4743 1783 4767
rect 41715 4801 41765 4825
rect 41715 4767 41723 4801
rect 41757 4767 41765 4801
rect 41715 4743 41765 4767
rect 1733 4465 1783 4489
rect 1733 4431 1741 4465
rect 1775 4431 1783 4465
rect 1733 4407 1783 4431
rect 41715 4465 41765 4489
rect 41715 4431 41723 4465
rect 41757 4431 41765 4465
rect 41715 4407 41765 4431
rect 1733 4129 1783 4153
rect 1733 4095 1741 4129
rect 1775 4095 1783 4129
rect 1733 4071 1783 4095
rect 41715 4129 41765 4153
rect 41715 4095 41723 4129
rect 41757 4095 41765 4129
rect 41715 4071 41765 4095
rect 1733 3793 1783 3817
rect 1733 3759 1741 3793
rect 1775 3759 1783 3793
rect 1733 3735 1783 3759
rect 41715 3793 41765 3817
rect 41715 3759 41723 3793
rect 41757 3759 41765 3793
rect 41715 3735 41765 3759
rect 1733 3457 1783 3481
rect 1733 3423 1741 3457
rect 1775 3423 1783 3457
rect 1733 3399 1783 3423
rect 41715 3457 41765 3481
rect 41715 3423 41723 3457
rect 41757 3423 41765 3457
rect 41715 3399 41765 3423
rect 1733 3121 1783 3145
rect 1733 3087 1741 3121
rect 1775 3087 1783 3121
rect 1733 3063 1783 3087
rect 41715 3121 41765 3145
rect 41715 3087 41723 3121
rect 41757 3087 41765 3121
rect 41715 3063 41765 3087
rect 1733 2785 1783 2809
rect 1733 2751 1741 2785
rect 1775 2751 1783 2785
rect 1733 2727 1783 2751
rect 41715 2785 41765 2809
rect 41715 2751 41723 2785
rect 41757 2751 41765 2785
rect 41715 2727 41765 2751
rect 1733 2449 1783 2473
rect 1733 2415 1741 2449
rect 1775 2415 1783 2449
rect 1733 2391 1783 2415
rect 41715 2449 41765 2473
rect 41715 2415 41723 2449
rect 41757 2415 41765 2449
rect 41715 2391 41765 2415
rect 1733 2113 1783 2137
rect 1733 2079 1741 2113
rect 1775 2079 1783 2113
rect 1733 2055 1783 2079
rect 41715 2113 41765 2137
rect 41715 2079 41723 2113
rect 41757 2079 41765 2113
rect 41715 2055 41765 2079
rect 2069 1777 2119 1801
rect 2069 1743 2077 1777
rect 2111 1743 2119 1777
rect 2069 1719 2119 1743
rect 2405 1777 2455 1801
rect 2405 1743 2413 1777
rect 2447 1743 2455 1777
rect 2405 1719 2455 1743
rect 2741 1777 2791 1801
rect 2741 1743 2749 1777
rect 2783 1743 2791 1777
rect 2741 1719 2791 1743
rect 3077 1777 3127 1801
rect 3077 1743 3085 1777
rect 3119 1743 3127 1777
rect 3077 1719 3127 1743
rect 3413 1777 3463 1801
rect 3413 1743 3421 1777
rect 3455 1743 3463 1777
rect 3413 1719 3463 1743
rect 3749 1777 3799 1801
rect 3749 1743 3757 1777
rect 3791 1743 3799 1777
rect 3749 1719 3799 1743
rect 4085 1777 4135 1801
rect 4085 1743 4093 1777
rect 4127 1743 4135 1777
rect 4085 1719 4135 1743
rect 4421 1777 4471 1801
rect 4421 1743 4429 1777
rect 4463 1743 4471 1777
rect 4421 1719 4471 1743
rect 4757 1777 4807 1801
rect 4757 1743 4765 1777
rect 4799 1743 4807 1777
rect 4757 1719 4807 1743
rect 5093 1777 5143 1801
rect 5093 1743 5101 1777
rect 5135 1743 5143 1777
rect 5093 1719 5143 1743
rect 5429 1777 5479 1801
rect 5429 1743 5437 1777
rect 5471 1743 5479 1777
rect 5429 1719 5479 1743
rect 5765 1777 5815 1801
rect 5765 1743 5773 1777
rect 5807 1743 5815 1777
rect 5765 1719 5815 1743
rect 6101 1777 6151 1801
rect 6101 1743 6109 1777
rect 6143 1743 6151 1777
rect 6101 1719 6151 1743
rect 6437 1777 6487 1801
rect 6437 1743 6445 1777
rect 6479 1743 6487 1777
rect 6437 1719 6487 1743
rect 6773 1777 6823 1801
rect 6773 1743 6781 1777
rect 6815 1743 6823 1777
rect 6773 1719 6823 1743
rect 7109 1777 7159 1801
rect 7109 1743 7117 1777
rect 7151 1743 7159 1777
rect 7109 1719 7159 1743
rect 7445 1777 7495 1801
rect 7445 1743 7453 1777
rect 7487 1743 7495 1777
rect 7445 1719 7495 1743
rect 7781 1777 7831 1801
rect 7781 1743 7789 1777
rect 7823 1743 7831 1777
rect 7781 1719 7831 1743
rect 8117 1777 8167 1801
rect 8117 1743 8125 1777
rect 8159 1743 8167 1777
rect 8117 1719 8167 1743
rect 8453 1777 8503 1801
rect 8453 1743 8461 1777
rect 8495 1743 8503 1777
rect 8453 1719 8503 1743
rect 8789 1777 8839 1801
rect 8789 1743 8797 1777
rect 8831 1743 8839 1777
rect 8789 1719 8839 1743
rect 9125 1777 9175 1801
rect 9125 1743 9133 1777
rect 9167 1743 9175 1777
rect 9125 1719 9175 1743
rect 9461 1777 9511 1801
rect 9461 1743 9469 1777
rect 9503 1743 9511 1777
rect 9461 1719 9511 1743
rect 9797 1777 9847 1801
rect 9797 1743 9805 1777
rect 9839 1743 9847 1777
rect 9797 1719 9847 1743
rect 10133 1777 10183 1801
rect 10133 1743 10141 1777
rect 10175 1743 10183 1777
rect 10133 1719 10183 1743
rect 10469 1777 10519 1801
rect 10469 1743 10477 1777
rect 10511 1743 10519 1777
rect 10469 1719 10519 1743
rect 10805 1777 10855 1801
rect 10805 1743 10813 1777
rect 10847 1743 10855 1777
rect 10805 1719 10855 1743
rect 11141 1777 11191 1801
rect 11141 1743 11149 1777
rect 11183 1743 11191 1777
rect 11141 1719 11191 1743
rect 11477 1777 11527 1801
rect 11477 1743 11485 1777
rect 11519 1743 11527 1777
rect 11477 1719 11527 1743
rect 11813 1777 11863 1801
rect 11813 1743 11821 1777
rect 11855 1743 11863 1777
rect 11813 1719 11863 1743
rect 12149 1777 12199 1801
rect 12149 1743 12157 1777
rect 12191 1743 12199 1777
rect 12149 1719 12199 1743
rect 12485 1777 12535 1801
rect 12485 1743 12493 1777
rect 12527 1743 12535 1777
rect 12485 1719 12535 1743
rect 12821 1777 12871 1801
rect 12821 1743 12829 1777
rect 12863 1743 12871 1777
rect 12821 1719 12871 1743
rect 13157 1777 13207 1801
rect 13157 1743 13165 1777
rect 13199 1743 13207 1777
rect 13157 1719 13207 1743
rect 13493 1777 13543 1801
rect 13493 1743 13501 1777
rect 13535 1743 13543 1777
rect 13493 1719 13543 1743
rect 13829 1777 13879 1801
rect 13829 1743 13837 1777
rect 13871 1743 13879 1777
rect 13829 1719 13879 1743
rect 14165 1777 14215 1801
rect 14165 1743 14173 1777
rect 14207 1743 14215 1777
rect 14165 1719 14215 1743
rect 14501 1777 14551 1801
rect 14501 1743 14509 1777
rect 14543 1743 14551 1777
rect 14501 1719 14551 1743
rect 14837 1777 14887 1801
rect 14837 1743 14845 1777
rect 14879 1743 14887 1777
rect 14837 1719 14887 1743
rect 15173 1777 15223 1801
rect 15173 1743 15181 1777
rect 15215 1743 15223 1777
rect 15173 1719 15223 1743
rect 15509 1777 15559 1801
rect 15509 1743 15517 1777
rect 15551 1743 15559 1777
rect 15509 1719 15559 1743
rect 15845 1777 15895 1801
rect 15845 1743 15853 1777
rect 15887 1743 15895 1777
rect 15845 1719 15895 1743
rect 16181 1777 16231 1801
rect 16181 1743 16189 1777
rect 16223 1743 16231 1777
rect 16181 1719 16231 1743
rect 16517 1777 16567 1801
rect 16517 1743 16525 1777
rect 16559 1743 16567 1777
rect 16517 1719 16567 1743
rect 16853 1777 16903 1801
rect 16853 1743 16861 1777
rect 16895 1743 16903 1777
rect 16853 1719 16903 1743
rect 17189 1777 17239 1801
rect 17189 1743 17197 1777
rect 17231 1743 17239 1777
rect 17189 1719 17239 1743
rect 17525 1777 17575 1801
rect 17525 1743 17533 1777
rect 17567 1743 17575 1777
rect 17525 1719 17575 1743
rect 17861 1777 17911 1801
rect 17861 1743 17869 1777
rect 17903 1743 17911 1777
rect 17861 1719 17911 1743
rect 18197 1777 18247 1801
rect 18197 1743 18205 1777
rect 18239 1743 18247 1777
rect 18197 1719 18247 1743
rect 18533 1777 18583 1801
rect 18533 1743 18541 1777
rect 18575 1743 18583 1777
rect 18533 1719 18583 1743
rect 18869 1777 18919 1801
rect 18869 1743 18877 1777
rect 18911 1743 18919 1777
rect 18869 1719 18919 1743
rect 19205 1777 19255 1801
rect 19205 1743 19213 1777
rect 19247 1743 19255 1777
rect 19205 1719 19255 1743
rect 19541 1777 19591 1801
rect 19541 1743 19549 1777
rect 19583 1743 19591 1777
rect 19541 1719 19591 1743
rect 19877 1777 19927 1801
rect 19877 1743 19885 1777
rect 19919 1743 19927 1777
rect 19877 1719 19927 1743
rect 20213 1777 20263 1801
rect 20213 1743 20221 1777
rect 20255 1743 20263 1777
rect 20213 1719 20263 1743
rect 20549 1777 20599 1801
rect 20549 1743 20557 1777
rect 20591 1743 20599 1777
rect 20549 1719 20599 1743
rect 20885 1777 20935 1801
rect 20885 1743 20893 1777
rect 20927 1743 20935 1777
rect 20885 1719 20935 1743
rect 21221 1777 21271 1801
rect 21221 1743 21229 1777
rect 21263 1743 21271 1777
rect 21221 1719 21271 1743
rect 21557 1777 21607 1801
rect 21557 1743 21565 1777
rect 21599 1743 21607 1777
rect 21557 1719 21607 1743
rect 21893 1777 21943 1801
rect 21893 1743 21901 1777
rect 21935 1743 21943 1777
rect 21893 1719 21943 1743
rect 22229 1777 22279 1801
rect 22229 1743 22237 1777
rect 22271 1743 22279 1777
rect 22229 1719 22279 1743
rect 22565 1777 22615 1801
rect 22565 1743 22573 1777
rect 22607 1743 22615 1777
rect 22565 1719 22615 1743
rect 22901 1777 22951 1801
rect 22901 1743 22909 1777
rect 22943 1743 22951 1777
rect 22901 1719 22951 1743
rect 23237 1777 23287 1801
rect 23237 1743 23245 1777
rect 23279 1743 23287 1777
rect 23237 1719 23287 1743
rect 23573 1777 23623 1801
rect 23573 1743 23581 1777
rect 23615 1743 23623 1777
rect 23573 1719 23623 1743
rect 23909 1777 23959 1801
rect 23909 1743 23917 1777
rect 23951 1743 23959 1777
rect 23909 1719 23959 1743
rect 24245 1777 24295 1801
rect 24245 1743 24253 1777
rect 24287 1743 24295 1777
rect 24245 1719 24295 1743
rect 24581 1777 24631 1801
rect 24581 1743 24589 1777
rect 24623 1743 24631 1777
rect 24581 1719 24631 1743
rect 24917 1777 24967 1801
rect 24917 1743 24925 1777
rect 24959 1743 24967 1777
rect 24917 1719 24967 1743
rect 25253 1777 25303 1801
rect 25253 1743 25261 1777
rect 25295 1743 25303 1777
rect 25253 1719 25303 1743
rect 25589 1777 25639 1801
rect 25589 1743 25597 1777
rect 25631 1743 25639 1777
rect 25589 1719 25639 1743
rect 25925 1777 25975 1801
rect 25925 1743 25933 1777
rect 25967 1743 25975 1777
rect 25925 1719 25975 1743
rect 26261 1777 26311 1801
rect 26261 1743 26269 1777
rect 26303 1743 26311 1777
rect 26261 1719 26311 1743
rect 26597 1777 26647 1801
rect 26597 1743 26605 1777
rect 26639 1743 26647 1777
rect 26597 1719 26647 1743
rect 26933 1777 26983 1801
rect 26933 1743 26941 1777
rect 26975 1743 26983 1777
rect 26933 1719 26983 1743
rect 27269 1777 27319 1801
rect 27269 1743 27277 1777
rect 27311 1743 27319 1777
rect 27269 1719 27319 1743
rect 27605 1777 27655 1801
rect 27605 1743 27613 1777
rect 27647 1743 27655 1777
rect 27605 1719 27655 1743
rect 27941 1777 27991 1801
rect 27941 1743 27949 1777
rect 27983 1743 27991 1777
rect 27941 1719 27991 1743
rect 28277 1777 28327 1801
rect 28277 1743 28285 1777
rect 28319 1743 28327 1777
rect 28277 1719 28327 1743
rect 28613 1777 28663 1801
rect 28613 1743 28621 1777
rect 28655 1743 28663 1777
rect 28613 1719 28663 1743
rect 28949 1777 28999 1801
rect 28949 1743 28957 1777
rect 28991 1743 28999 1777
rect 28949 1719 28999 1743
rect 29285 1777 29335 1801
rect 29285 1743 29293 1777
rect 29327 1743 29335 1777
rect 29285 1719 29335 1743
rect 29621 1777 29671 1801
rect 29621 1743 29629 1777
rect 29663 1743 29671 1777
rect 29621 1719 29671 1743
rect 29957 1777 30007 1801
rect 29957 1743 29965 1777
rect 29999 1743 30007 1777
rect 29957 1719 30007 1743
rect 30293 1777 30343 1801
rect 30293 1743 30301 1777
rect 30335 1743 30343 1777
rect 30293 1719 30343 1743
rect 30629 1777 30679 1801
rect 30629 1743 30637 1777
rect 30671 1743 30679 1777
rect 30629 1719 30679 1743
rect 30965 1777 31015 1801
rect 30965 1743 30973 1777
rect 31007 1743 31015 1777
rect 30965 1719 31015 1743
rect 31301 1777 31351 1801
rect 31301 1743 31309 1777
rect 31343 1743 31351 1777
rect 31301 1719 31351 1743
rect 31637 1777 31687 1801
rect 31637 1743 31645 1777
rect 31679 1743 31687 1777
rect 31637 1719 31687 1743
rect 31973 1777 32023 1801
rect 31973 1743 31981 1777
rect 32015 1743 32023 1777
rect 31973 1719 32023 1743
rect 32309 1777 32359 1801
rect 32309 1743 32317 1777
rect 32351 1743 32359 1777
rect 32309 1719 32359 1743
rect 32645 1777 32695 1801
rect 32645 1743 32653 1777
rect 32687 1743 32695 1777
rect 32645 1719 32695 1743
rect 32981 1777 33031 1801
rect 32981 1743 32989 1777
rect 33023 1743 33031 1777
rect 32981 1719 33031 1743
rect 33317 1777 33367 1801
rect 33317 1743 33325 1777
rect 33359 1743 33367 1777
rect 33317 1719 33367 1743
rect 33653 1777 33703 1801
rect 33653 1743 33661 1777
rect 33695 1743 33703 1777
rect 33653 1719 33703 1743
rect 33989 1777 34039 1801
rect 33989 1743 33997 1777
rect 34031 1743 34039 1777
rect 33989 1719 34039 1743
rect 34325 1777 34375 1801
rect 34325 1743 34333 1777
rect 34367 1743 34375 1777
rect 34325 1719 34375 1743
rect 34661 1777 34711 1801
rect 34661 1743 34669 1777
rect 34703 1743 34711 1777
rect 34661 1719 34711 1743
rect 34997 1777 35047 1801
rect 34997 1743 35005 1777
rect 35039 1743 35047 1777
rect 34997 1719 35047 1743
rect 35333 1777 35383 1801
rect 35333 1743 35341 1777
rect 35375 1743 35383 1777
rect 35333 1719 35383 1743
rect 35669 1777 35719 1801
rect 35669 1743 35677 1777
rect 35711 1743 35719 1777
rect 35669 1719 35719 1743
rect 36005 1777 36055 1801
rect 36005 1743 36013 1777
rect 36047 1743 36055 1777
rect 36005 1719 36055 1743
rect 36341 1777 36391 1801
rect 36341 1743 36349 1777
rect 36383 1743 36391 1777
rect 36341 1719 36391 1743
rect 36677 1777 36727 1801
rect 36677 1743 36685 1777
rect 36719 1743 36727 1777
rect 36677 1719 36727 1743
rect 37013 1777 37063 1801
rect 37013 1743 37021 1777
rect 37055 1743 37063 1777
rect 37013 1719 37063 1743
rect 37349 1777 37399 1801
rect 37349 1743 37357 1777
rect 37391 1743 37399 1777
rect 37349 1719 37399 1743
rect 37685 1777 37735 1801
rect 37685 1743 37693 1777
rect 37727 1743 37735 1777
rect 37685 1719 37735 1743
rect 38021 1777 38071 1801
rect 38021 1743 38029 1777
rect 38063 1743 38071 1777
rect 38021 1719 38071 1743
rect 38357 1777 38407 1801
rect 38357 1743 38365 1777
rect 38399 1743 38407 1777
rect 38357 1719 38407 1743
rect 38693 1777 38743 1801
rect 38693 1743 38701 1777
rect 38735 1743 38743 1777
rect 38693 1719 38743 1743
rect 39029 1777 39079 1801
rect 39029 1743 39037 1777
rect 39071 1743 39079 1777
rect 39029 1719 39079 1743
rect 39365 1777 39415 1801
rect 39365 1743 39373 1777
rect 39407 1743 39415 1777
rect 39365 1719 39415 1743
rect 39701 1777 39751 1801
rect 39701 1743 39709 1777
rect 39743 1743 39751 1777
rect 39701 1719 39751 1743
rect 40037 1777 40087 1801
rect 40037 1743 40045 1777
rect 40079 1743 40087 1777
rect 40037 1719 40087 1743
rect 40373 1777 40423 1801
rect 40373 1743 40381 1777
rect 40415 1743 40423 1777
rect 40373 1719 40423 1743
rect 40709 1777 40759 1801
rect 40709 1743 40717 1777
rect 40751 1743 40759 1777
rect 40709 1719 40759 1743
rect 41045 1777 41095 1801
rect 41045 1743 41053 1777
rect 41087 1743 41095 1777
rect 41045 1719 41095 1743
<< nsubdiffcont >>
rect 2077 31367 2111 31401
rect 2413 31367 2447 31401
rect 2749 31367 2783 31401
rect 3085 31367 3119 31401
rect 3421 31367 3455 31401
rect 3757 31367 3791 31401
rect 4093 31367 4127 31401
rect 4429 31367 4463 31401
rect 4765 31367 4799 31401
rect 5101 31367 5135 31401
rect 5437 31367 5471 31401
rect 5773 31367 5807 31401
rect 6109 31367 6143 31401
rect 6445 31367 6479 31401
rect 6781 31367 6815 31401
rect 7117 31367 7151 31401
rect 7453 31367 7487 31401
rect 7789 31367 7823 31401
rect 8125 31367 8159 31401
rect 8461 31367 8495 31401
rect 8797 31367 8831 31401
rect 9133 31367 9167 31401
rect 9469 31367 9503 31401
rect 9805 31367 9839 31401
rect 10141 31367 10175 31401
rect 10477 31367 10511 31401
rect 10813 31367 10847 31401
rect 11149 31367 11183 31401
rect 11485 31367 11519 31401
rect 11821 31367 11855 31401
rect 12157 31367 12191 31401
rect 12493 31367 12527 31401
rect 12829 31367 12863 31401
rect 13165 31367 13199 31401
rect 13501 31367 13535 31401
rect 13837 31367 13871 31401
rect 14173 31367 14207 31401
rect 14509 31367 14543 31401
rect 14845 31367 14879 31401
rect 15181 31367 15215 31401
rect 15517 31367 15551 31401
rect 15853 31367 15887 31401
rect 16189 31367 16223 31401
rect 16525 31367 16559 31401
rect 16861 31367 16895 31401
rect 17197 31367 17231 31401
rect 17533 31367 17567 31401
rect 17869 31367 17903 31401
rect 18205 31367 18239 31401
rect 18541 31367 18575 31401
rect 18877 31367 18911 31401
rect 19213 31367 19247 31401
rect 19549 31367 19583 31401
rect 19885 31367 19919 31401
rect 20221 31367 20255 31401
rect 20557 31367 20591 31401
rect 20893 31367 20927 31401
rect 21229 31367 21263 31401
rect 21565 31367 21599 31401
rect 21901 31367 21935 31401
rect 22237 31367 22271 31401
rect 22573 31367 22607 31401
rect 22909 31367 22943 31401
rect 23245 31367 23279 31401
rect 23581 31367 23615 31401
rect 23917 31367 23951 31401
rect 24253 31367 24287 31401
rect 24589 31367 24623 31401
rect 24925 31367 24959 31401
rect 25261 31367 25295 31401
rect 25597 31367 25631 31401
rect 25933 31367 25967 31401
rect 26269 31367 26303 31401
rect 26605 31367 26639 31401
rect 26941 31367 26975 31401
rect 27277 31367 27311 31401
rect 27613 31367 27647 31401
rect 27949 31367 27983 31401
rect 28285 31367 28319 31401
rect 28621 31367 28655 31401
rect 28957 31367 28991 31401
rect 29293 31367 29327 31401
rect 29629 31367 29663 31401
rect 29965 31367 29999 31401
rect 30301 31367 30335 31401
rect 30637 31367 30671 31401
rect 30973 31367 31007 31401
rect 31309 31367 31343 31401
rect 31645 31367 31679 31401
rect 31981 31367 32015 31401
rect 32317 31367 32351 31401
rect 32653 31367 32687 31401
rect 32989 31367 33023 31401
rect 33325 31367 33359 31401
rect 33661 31367 33695 31401
rect 33997 31367 34031 31401
rect 34333 31367 34367 31401
rect 34669 31367 34703 31401
rect 35005 31367 35039 31401
rect 35341 31367 35375 31401
rect 35677 31367 35711 31401
rect 36013 31367 36047 31401
rect 36349 31367 36383 31401
rect 36685 31367 36719 31401
rect 37021 31367 37055 31401
rect 37357 31367 37391 31401
rect 37693 31367 37727 31401
rect 38029 31367 38063 31401
rect 38365 31367 38399 31401
rect 38701 31367 38735 31401
rect 39037 31367 39071 31401
rect 39373 31367 39407 31401
rect 39709 31367 39743 31401
rect 40045 31367 40079 31401
rect 40381 31367 40415 31401
rect 40717 31367 40751 31401
rect 41053 31367 41087 31401
rect 1741 30975 1775 31009
rect 41723 30975 41757 31009
rect 1741 30639 1775 30673
rect 41723 30639 41757 30673
rect 1741 30303 1775 30337
rect 41723 30303 41757 30337
rect 1741 29967 1775 30001
rect 41723 29967 41757 30001
rect 1741 29631 1775 29665
rect 41723 29631 41757 29665
rect 1741 29295 1775 29329
rect 41723 29295 41757 29329
rect 1741 28959 1775 28993
rect 41723 28959 41757 28993
rect 1741 28623 1775 28657
rect 41723 28623 41757 28657
rect 1741 28287 1775 28321
rect 41723 28287 41757 28321
rect 1741 27951 1775 27985
rect 41723 27951 41757 27985
rect 1741 27615 1775 27649
rect 41723 27615 41757 27649
rect 1741 27279 1775 27313
rect 41723 27279 41757 27313
rect 1741 26943 1775 26977
rect 41723 26943 41757 26977
rect 1741 26607 1775 26641
rect 41723 26607 41757 26641
rect 1741 26271 1775 26305
rect 41723 26271 41757 26305
rect 1741 25935 1775 25969
rect 41723 25935 41757 25969
rect 1741 25599 1775 25633
rect 41723 25599 41757 25633
rect 1741 25263 1775 25297
rect 41723 25263 41757 25297
rect 1741 24927 1775 24961
rect 41723 24927 41757 24961
rect 1741 24591 1775 24625
rect 41723 24591 41757 24625
rect 1741 24255 1775 24289
rect 41723 24255 41757 24289
rect 1741 23919 1775 23953
rect 41723 23919 41757 23953
rect 1741 23583 1775 23617
rect 41723 23583 41757 23617
rect 1741 23247 1775 23281
rect 41723 23247 41757 23281
rect 1741 22911 1775 22945
rect 41723 22911 41757 22945
rect 1741 22575 1775 22609
rect 41723 22575 41757 22609
rect 1741 22239 1775 22273
rect 41723 22239 41757 22273
rect 1741 21903 1775 21937
rect 41723 21903 41757 21937
rect 1741 21567 1775 21601
rect 41723 21567 41757 21601
rect 1741 21231 1775 21265
rect 41723 21231 41757 21265
rect 1741 20895 1775 20929
rect 41723 20895 41757 20929
rect 1741 20559 1775 20593
rect 41723 20559 41757 20593
rect 1741 20223 1775 20257
rect 41723 20223 41757 20257
rect 1741 19887 1775 19921
rect 41723 19887 41757 19921
rect 1741 19551 1775 19585
rect 41723 19551 41757 19585
rect 1741 19215 1775 19249
rect 41723 19215 41757 19249
rect 1741 18879 1775 18913
rect 41723 18879 41757 18913
rect 1741 18543 1775 18577
rect 41723 18543 41757 18577
rect 1741 18207 1775 18241
rect 41723 18207 41757 18241
rect 1741 17871 1775 17905
rect 41723 17871 41757 17905
rect 1741 17535 1775 17569
rect 41723 17535 41757 17569
rect 1741 17199 1775 17233
rect 41723 17199 41757 17233
rect 1741 16863 1775 16897
rect 41723 16863 41757 16897
rect 1741 16527 1775 16561
rect 41723 16527 41757 16561
rect 1741 16191 1775 16225
rect 41723 16191 41757 16225
rect 1741 15855 1775 15889
rect 41723 15855 41757 15889
rect 1741 15519 1775 15553
rect 41723 15519 41757 15553
rect 1741 15183 1775 15217
rect 41723 15183 41757 15217
rect 1741 14847 1775 14881
rect 41723 14847 41757 14881
rect 1741 14511 1775 14545
rect 41723 14511 41757 14545
rect 1741 14175 1775 14209
rect 41723 14175 41757 14209
rect 1741 13839 1775 13873
rect 41723 13839 41757 13873
rect 1741 13503 1775 13537
rect 41723 13503 41757 13537
rect 1741 13167 1775 13201
rect 41723 13167 41757 13201
rect 1741 12831 1775 12865
rect 41723 12831 41757 12865
rect 1741 12495 1775 12529
rect 41723 12495 41757 12529
rect 1741 12159 1775 12193
rect 41723 12159 41757 12193
rect 1741 11823 1775 11857
rect 41723 11823 41757 11857
rect 1741 11487 1775 11521
rect 41723 11487 41757 11521
rect 1741 11151 1775 11185
rect 41723 11151 41757 11185
rect 1741 10815 1775 10849
rect 41723 10815 41757 10849
rect 1741 10479 1775 10513
rect 41723 10479 41757 10513
rect 1741 10143 1775 10177
rect 41723 10143 41757 10177
rect 1741 9807 1775 9841
rect 41723 9807 41757 9841
rect 1741 9471 1775 9505
rect 41723 9471 41757 9505
rect 1741 9135 1775 9169
rect 41723 9135 41757 9169
rect 1741 8799 1775 8833
rect 41723 8799 41757 8833
rect 1741 8463 1775 8497
rect 41723 8463 41757 8497
rect 1741 8127 1775 8161
rect 41723 8127 41757 8161
rect 1741 7791 1775 7825
rect 41723 7791 41757 7825
rect 1741 7455 1775 7489
rect 41723 7455 41757 7489
rect 1741 7119 1775 7153
rect 41723 7119 41757 7153
rect 1741 6783 1775 6817
rect 41723 6783 41757 6817
rect 1741 6447 1775 6481
rect 41723 6447 41757 6481
rect 1741 6111 1775 6145
rect 41723 6111 41757 6145
rect 1741 5775 1775 5809
rect 41723 5775 41757 5809
rect 1741 5439 1775 5473
rect 41723 5439 41757 5473
rect 1741 5103 1775 5137
rect 41723 5103 41757 5137
rect 1741 4767 1775 4801
rect 41723 4767 41757 4801
rect 1741 4431 1775 4465
rect 41723 4431 41757 4465
rect 1741 4095 1775 4129
rect 41723 4095 41757 4129
rect 1741 3759 1775 3793
rect 41723 3759 41757 3793
rect 1741 3423 1775 3457
rect 41723 3423 41757 3457
rect 1741 3087 1775 3121
rect 41723 3087 41757 3121
rect 1741 2751 1775 2785
rect 41723 2751 41757 2785
rect 1741 2415 1775 2449
rect 41723 2415 41757 2449
rect 1741 2079 1775 2113
rect 41723 2079 41757 2113
rect 2077 1743 2111 1777
rect 2413 1743 2447 1777
rect 2749 1743 2783 1777
rect 3085 1743 3119 1777
rect 3421 1743 3455 1777
rect 3757 1743 3791 1777
rect 4093 1743 4127 1777
rect 4429 1743 4463 1777
rect 4765 1743 4799 1777
rect 5101 1743 5135 1777
rect 5437 1743 5471 1777
rect 5773 1743 5807 1777
rect 6109 1743 6143 1777
rect 6445 1743 6479 1777
rect 6781 1743 6815 1777
rect 7117 1743 7151 1777
rect 7453 1743 7487 1777
rect 7789 1743 7823 1777
rect 8125 1743 8159 1777
rect 8461 1743 8495 1777
rect 8797 1743 8831 1777
rect 9133 1743 9167 1777
rect 9469 1743 9503 1777
rect 9805 1743 9839 1777
rect 10141 1743 10175 1777
rect 10477 1743 10511 1777
rect 10813 1743 10847 1777
rect 11149 1743 11183 1777
rect 11485 1743 11519 1777
rect 11821 1743 11855 1777
rect 12157 1743 12191 1777
rect 12493 1743 12527 1777
rect 12829 1743 12863 1777
rect 13165 1743 13199 1777
rect 13501 1743 13535 1777
rect 13837 1743 13871 1777
rect 14173 1743 14207 1777
rect 14509 1743 14543 1777
rect 14845 1743 14879 1777
rect 15181 1743 15215 1777
rect 15517 1743 15551 1777
rect 15853 1743 15887 1777
rect 16189 1743 16223 1777
rect 16525 1743 16559 1777
rect 16861 1743 16895 1777
rect 17197 1743 17231 1777
rect 17533 1743 17567 1777
rect 17869 1743 17903 1777
rect 18205 1743 18239 1777
rect 18541 1743 18575 1777
rect 18877 1743 18911 1777
rect 19213 1743 19247 1777
rect 19549 1743 19583 1777
rect 19885 1743 19919 1777
rect 20221 1743 20255 1777
rect 20557 1743 20591 1777
rect 20893 1743 20927 1777
rect 21229 1743 21263 1777
rect 21565 1743 21599 1777
rect 21901 1743 21935 1777
rect 22237 1743 22271 1777
rect 22573 1743 22607 1777
rect 22909 1743 22943 1777
rect 23245 1743 23279 1777
rect 23581 1743 23615 1777
rect 23917 1743 23951 1777
rect 24253 1743 24287 1777
rect 24589 1743 24623 1777
rect 24925 1743 24959 1777
rect 25261 1743 25295 1777
rect 25597 1743 25631 1777
rect 25933 1743 25967 1777
rect 26269 1743 26303 1777
rect 26605 1743 26639 1777
rect 26941 1743 26975 1777
rect 27277 1743 27311 1777
rect 27613 1743 27647 1777
rect 27949 1743 27983 1777
rect 28285 1743 28319 1777
rect 28621 1743 28655 1777
rect 28957 1743 28991 1777
rect 29293 1743 29327 1777
rect 29629 1743 29663 1777
rect 29965 1743 29999 1777
rect 30301 1743 30335 1777
rect 30637 1743 30671 1777
rect 30973 1743 31007 1777
rect 31309 1743 31343 1777
rect 31645 1743 31679 1777
rect 31981 1743 32015 1777
rect 32317 1743 32351 1777
rect 32653 1743 32687 1777
rect 32989 1743 33023 1777
rect 33325 1743 33359 1777
rect 33661 1743 33695 1777
rect 33997 1743 34031 1777
rect 34333 1743 34367 1777
rect 34669 1743 34703 1777
rect 35005 1743 35039 1777
rect 35341 1743 35375 1777
rect 35677 1743 35711 1777
rect 36013 1743 36047 1777
rect 36349 1743 36383 1777
rect 36685 1743 36719 1777
rect 37021 1743 37055 1777
rect 37357 1743 37391 1777
rect 37693 1743 37727 1777
rect 38029 1743 38063 1777
rect 38365 1743 38399 1777
rect 38701 1743 38735 1777
rect 39037 1743 39071 1777
rect 39373 1743 39407 1777
rect 39709 1743 39743 1777
rect 40045 1743 40079 1777
rect 40381 1743 40415 1777
rect 40717 1743 40751 1777
rect 41053 1743 41087 1777
<< locali >>
rect 2077 31401 2111 31417
rect 2077 31351 2111 31367
rect 2413 31401 2447 31417
rect 2413 31351 2447 31367
rect 2749 31401 2783 31417
rect 2749 31351 2783 31367
rect 3085 31401 3119 31417
rect 3085 31351 3119 31367
rect 3421 31401 3455 31417
rect 3421 31351 3455 31367
rect 3757 31401 3791 31417
rect 3757 31351 3791 31367
rect 4093 31401 4127 31417
rect 4093 31351 4127 31367
rect 4429 31401 4463 31417
rect 4429 31351 4463 31367
rect 4765 31401 4799 31417
rect 4765 31351 4799 31367
rect 5101 31401 5135 31417
rect 5101 31351 5135 31367
rect 5437 31401 5471 31417
rect 5437 31351 5471 31367
rect 5773 31401 5807 31417
rect 5773 31351 5807 31367
rect 6109 31401 6143 31417
rect 6109 31351 6143 31367
rect 6445 31401 6479 31417
rect 6445 31351 6479 31367
rect 6781 31401 6815 31417
rect 6781 31351 6815 31367
rect 7117 31401 7151 31417
rect 7117 31351 7151 31367
rect 7453 31401 7487 31417
rect 7453 31351 7487 31367
rect 7789 31401 7823 31417
rect 7789 31351 7823 31367
rect 8125 31401 8159 31417
rect 8125 31351 8159 31367
rect 8461 31401 8495 31417
rect 8461 31351 8495 31367
rect 8797 31401 8831 31417
rect 8797 31351 8831 31367
rect 9133 31401 9167 31417
rect 9133 31351 9167 31367
rect 9469 31401 9503 31417
rect 9469 31351 9503 31367
rect 9805 31401 9839 31417
rect 9805 31351 9839 31367
rect 10141 31401 10175 31417
rect 10141 31351 10175 31367
rect 10477 31401 10511 31417
rect 10477 31351 10511 31367
rect 10813 31401 10847 31417
rect 10813 31351 10847 31367
rect 11149 31401 11183 31417
rect 11149 31351 11183 31367
rect 11485 31401 11519 31417
rect 11485 31351 11519 31367
rect 11821 31401 11855 31417
rect 11821 31351 11855 31367
rect 12157 31401 12191 31417
rect 12157 31351 12191 31367
rect 12493 31401 12527 31417
rect 12493 31351 12527 31367
rect 12829 31401 12863 31417
rect 12829 31351 12863 31367
rect 13165 31401 13199 31417
rect 13165 31351 13199 31367
rect 13501 31401 13535 31417
rect 13501 31351 13535 31367
rect 13837 31401 13871 31417
rect 13837 31351 13871 31367
rect 14173 31401 14207 31417
rect 14173 31351 14207 31367
rect 14509 31401 14543 31417
rect 14509 31351 14543 31367
rect 14845 31401 14879 31417
rect 14845 31351 14879 31367
rect 15181 31401 15215 31417
rect 15181 31351 15215 31367
rect 15517 31401 15551 31417
rect 15517 31351 15551 31367
rect 15853 31401 15887 31417
rect 15853 31351 15887 31367
rect 16189 31401 16223 31417
rect 16189 31351 16223 31367
rect 16525 31401 16559 31417
rect 16525 31351 16559 31367
rect 16861 31401 16895 31417
rect 16861 31351 16895 31367
rect 17197 31401 17231 31417
rect 17197 31351 17231 31367
rect 17533 31401 17567 31417
rect 17533 31351 17567 31367
rect 17869 31401 17903 31417
rect 17869 31351 17903 31367
rect 18205 31401 18239 31417
rect 18205 31351 18239 31367
rect 18541 31401 18575 31417
rect 18541 31351 18575 31367
rect 18877 31401 18911 31417
rect 18877 31351 18911 31367
rect 19213 31401 19247 31417
rect 19213 31351 19247 31367
rect 19549 31401 19583 31417
rect 19549 31351 19583 31367
rect 19885 31401 19919 31417
rect 19885 31351 19919 31367
rect 20221 31401 20255 31417
rect 20221 31351 20255 31367
rect 20557 31401 20591 31417
rect 20557 31351 20591 31367
rect 20893 31401 20927 31417
rect 20893 31351 20927 31367
rect 21229 31401 21263 31417
rect 21229 31351 21263 31367
rect 21565 31401 21599 31417
rect 21565 31351 21599 31367
rect 21901 31401 21935 31417
rect 21901 31351 21935 31367
rect 22237 31401 22271 31417
rect 22237 31351 22271 31367
rect 22573 31401 22607 31417
rect 22573 31351 22607 31367
rect 22909 31401 22943 31417
rect 22909 31351 22943 31367
rect 23245 31401 23279 31417
rect 23245 31351 23279 31367
rect 23581 31401 23615 31417
rect 23581 31351 23615 31367
rect 23917 31401 23951 31417
rect 23917 31351 23951 31367
rect 24253 31401 24287 31417
rect 24253 31351 24287 31367
rect 24589 31401 24623 31417
rect 24589 31351 24623 31367
rect 24925 31401 24959 31417
rect 24925 31351 24959 31367
rect 25261 31401 25295 31417
rect 25261 31351 25295 31367
rect 25597 31401 25631 31417
rect 25597 31351 25631 31367
rect 25933 31401 25967 31417
rect 25933 31351 25967 31367
rect 26269 31401 26303 31417
rect 26269 31351 26303 31367
rect 26605 31401 26639 31417
rect 26605 31351 26639 31367
rect 26941 31401 26975 31417
rect 26941 31351 26975 31367
rect 27277 31401 27311 31417
rect 27277 31351 27311 31367
rect 27613 31401 27647 31417
rect 27613 31351 27647 31367
rect 27949 31401 27983 31417
rect 27949 31351 27983 31367
rect 28285 31401 28319 31417
rect 28285 31351 28319 31367
rect 28621 31401 28655 31417
rect 28621 31351 28655 31367
rect 28957 31401 28991 31417
rect 28957 31351 28991 31367
rect 29293 31401 29327 31417
rect 29293 31351 29327 31367
rect 29629 31401 29663 31417
rect 29629 31351 29663 31367
rect 29965 31401 29999 31417
rect 29965 31351 29999 31367
rect 30301 31401 30335 31417
rect 30301 31351 30335 31367
rect 30637 31401 30671 31417
rect 30637 31351 30671 31367
rect 30973 31401 31007 31417
rect 30973 31351 31007 31367
rect 31309 31401 31343 31417
rect 31309 31351 31343 31367
rect 31645 31401 31679 31417
rect 31645 31351 31679 31367
rect 31981 31401 32015 31417
rect 31981 31351 32015 31367
rect 32317 31401 32351 31417
rect 32317 31351 32351 31367
rect 32653 31401 32687 31417
rect 32653 31351 32687 31367
rect 32989 31401 33023 31417
rect 32989 31351 33023 31367
rect 33325 31401 33359 31417
rect 33325 31351 33359 31367
rect 33661 31401 33695 31417
rect 33661 31351 33695 31367
rect 33997 31401 34031 31417
rect 33997 31351 34031 31367
rect 34333 31401 34367 31417
rect 34333 31351 34367 31367
rect 34669 31401 34703 31417
rect 34669 31351 34703 31367
rect 35005 31401 35039 31417
rect 35005 31351 35039 31367
rect 35341 31401 35375 31417
rect 35341 31351 35375 31367
rect 35677 31401 35711 31417
rect 35677 31351 35711 31367
rect 36013 31401 36047 31417
rect 36013 31351 36047 31367
rect 36349 31401 36383 31417
rect 36349 31351 36383 31367
rect 36685 31401 36719 31417
rect 36685 31351 36719 31367
rect 37021 31401 37055 31417
rect 37021 31351 37055 31367
rect 37357 31401 37391 31417
rect 37357 31351 37391 31367
rect 37693 31401 37727 31417
rect 37693 31351 37727 31367
rect 38029 31401 38063 31417
rect 38029 31351 38063 31367
rect 38365 31401 38399 31417
rect 38365 31351 38399 31367
rect 38701 31401 38735 31417
rect 38701 31351 38735 31367
rect 39037 31401 39071 31417
rect 39037 31351 39071 31367
rect 39373 31401 39407 31417
rect 39373 31351 39407 31367
rect 39709 31401 39743 31417
rect 39709 31351 39743 31367
rect 40045 31401 40079 31417
rect 40045 31351 40079 31367
rect 40381 31401 40415 31417
rect 40381 31351 40415 31367
rect 40717 31401 40751 31417
rect 40717 31351 40751 31367
rect 41053 31401 41087 31417
rect 41053 31351 41087 31367
rect 1741 31009 1775 31025
rect 1741 30959 1775 30975
rect 41723 31009 41757 31025
rect 41723 30959 41757 30975
rect 1741 30673 1775 30689
rect 1741 30623 1775 30639
rect 41723 30673 41757 30689
rect 41723 30623 41757 30639
rect 1741 30337 1775 30353
rect 1741 30287 1775 30303
rect 41723 30337 41757 30353
rect 41723 30287 41757 30303
rect 1741 30001 1775 30017
rect 1741 29951 1775 29967
rect 41723 30001 41757 30017
rect 41723 29951 41757 29967
rect 1741 29665 1775 29681
rect 1741 29615 1775 29631
rect 41723 29665 41757 29681
rect 41723 29615 41757 29631
rect 1741 29329 1775 29345
rect 1741 29279 1775 29295
rect 41723 29329 41757 29345
rect 41723 29279 41757 29295
rect 1741 28993 1775 29009
rect 1741 28943 1775 28959
rect 41723 28993 41757 29009
rect 41723 28943 41757 28959
rect 1741 28657 1775 28673
rect 1741 28607 1775 28623
rect 41723 28657 41757 28673
rect 41723 28607 41757 28623
rect 1741 28321 1775 28337
rect 1741 28271 1775 28287
rect 41723 28321 41757 28337
rect 41723 28271 41757 28287
rect 1741 27985 1775 28001
rect 1741 27935 1775 27951
rect 41723 27985 41757 28001
rect 41723 27935 41757 27951
rect 1741 27649 1775 27665
rect 1741 27599 1775 27615
rect 41723 27649 41757 27665
rect 41723 27599 41757 27615
rect 1741 27313 1775 27329
rect 1741 27263 1775 27279
rect 41723 27313 41757 27329
rect 41723 27263 41757 27279
rect 1741 26977 1775 26993
rect 1741 26927 1775 26943
rect 41723 26977 41757 26993
rect 41723 26927 41757 26943
rect 1741 26641 1775 26657
rect 1741 26591 1775 26607
rect 41723 26641 41757 26657
rect 41723 26591 41757 26607
rect 1741 26305 1775 26321
rect 1741 26255 1775 26271
rect 41723 26305 41757 26321
rect 41723 26255 41757 26271
rect 1741 25969 1775 25985
rect 1741 25919 1775 25935
rect 41723 25969 41757 25985
rect 41723 25919 41757 25935
rect 1741 25633 1775 25649
rect 1741 25583 1775 25599
rect 41723 25633 41757 25649
rect 41723 25583 41757 25599
rect 1741 25297 1775 25313
rect 1741 25247 1775 25263
rect 41723 25297 41757 25313
rect 41723 25247 41757 25263
rect 1741 24961 1775 24977
rect 1741 24911 1775 24927
rect 41723 24961 41757 24977
rect 41723 24911 41757 24927
rect 1741 24625 1775 24641
rect 1741 24575 1775 24591
rect 41723 24625 41757 24641
rect 41723 24575 41757 24591
rect 1741 24289 1775 24305
rect 1741 24239 1775 24255
rect 41723 24289 41757 24305
rect 41723 24239 41757 24255
rect 1741 23953 1775 23969
rect 1741 23903 1775 23919
rect 41723 23953 41757 23969
rect 41723 23903 41757 23919
rect 1741 23617 1775 23633
rect 1741 23567 1775 23583
rect 41723 23617 41757 23633
rect 41723 23567 41757 23583
rect 1741 23281 1775 23297
rect 1741 23231 1775 23247
rect 41723 23281 41757 23297
rect 41723 23231 41757 23247
rect 1741 22945 1775 22961
rect 1741 22895 1775 22911
rect 41723 22945 41757 22961
rect 41723 22895 41757 22911
rect 1741 22609 1775 22625
rect 1741 22559 1775 22575
rect 41723 22609 41757 22625
rect 41723 22559 41757 22575
rect 1741 22273 1775 22289
rect 1741 22223 1775 22239
rect 41723 22273 41757 22289
rect 41723 22223 41757 22239
rect 1741 21937 1775 21953
rect 1741 21887 1775 21903
rect 41723 21937 41757 21953
rect 41723 21887 41757 21903
rect 1741 21601 1775 21617
rect 1741 21551 1775 21567
rect 41723 21601 41757 21617
rect 41723 21551 41757 21567
rect 1741 21265 1775 21281
rect 1741 21215 1775 21231
rect 41723 21265 41757 21281
rect 41723 21215 41757 21231
rect 1741 20929 1775 20945
rect 1741 20879 1775 20895
rect 41723 20929 41757 20945
rect 41723 20879 41757 20895
rect 1741 20593 1775 20609
rect 1741 20543 1775 20559
rect 41723 20593 41757 20609
rect 41723 20543 41757 20559
rect 1741 20257 1775 20273
rect 1741 20207 1775 20223
rect 41723 20257 41757 20273
rect 41723 20207 41757 20223
rect 1741 19921 1775 19937
rect 1741 19871 1775 19887
rect 41723 19921 41757 19937
rect 41723 19871 41757 19887
rect 1741 19585 1775 19601
rect 1741 19535 1775 19551
rect 41723 19585 41757 19601
rect 41723 19535 41757 19551
rect 1741 19249 1775 19265
rect 1741 19199 1775 19215
rect 41723 19249 41757 19265
rect 41723 19199 41757 19215
rect 1741 18913 1775 18929
rect 1741 18863 1775 18879
rect 41723 18913 41757 18929
rect 41723 18863 41757 18879
rect 1741 18577 1775 18593
rect 1741 18527 1775 18543
rect 41723 18577 41757 18593
rect 41723 18527 41757 18543
rect 1741 18241 1775 18257
rect 1741 18191 1775 18207
rect 41723 18241 41757 18257
rect 41723 18191 41757 18207
rect 1741 17905 1775 17921
rect 1741 17855 1775 17871
rect 41723 17905 41757 17921
rect 41723 17855 41757 17871
rect 1741 17569 1775 17585
rect 1741 17519 1775 17535
rect 41723 17569 41757 17585
rect 41723 17519 41757 17535
rect 1741 17233 1775 17249
rect 1741 17183 1775 17199
rect 41723 17233 41757 17249
rect 41723 17183 41757 17199
rect 1741 16897 1775 16913
rect 1741 16847 1775 16863
rect 41723 16897 41757 16913
rect 41723 16847 41757 16863
rect 1741 16561 1775 16577
rect 1741 16511 1775 16527
rect 41723 16561 41757 16577
rect 41723 16511 41757 16527
rect 1741 16225 1775 16241
rect 1741 16175 1775 16191
rect 41723 16225 41757 16241
rect 41723 16175 41757 16191
rect 1741 15889 1775 15905
rect 1741 15839 1775 15855
rect 41723 15889 41757 15905
rect 41723 15839 41757 15855
rect 1741 15553 1775 15569
rect 1741 15503 1775 15519
rect 41723 15553 41757 15569
rect 41723 15503 41757 15519
rect 1741 15217 1775 15233
rect 1741 15167 1775 15183
rect 41723 15217 41757 15233
rect 41723 15167 41757 15183
rect 1741 14881 1775 14897
rect 1741 14831 1775 14847
rect 41723 14881 41757 14897
rect 41723 14831 41757 14847
rect 1741 14545 1775 14561
rect 1741 14495 1775 14511
rect 41723 14545 41757 14561
rect 41723 14495 41757 14511
rect 1741 14209 1775 14225
rect 1741 14159 1775 14175
rect 41723 14209 41757 14225
rect 41723 14159 41757 14175
rect 1741 13873 1775 13889
rect 1741 13823 1775 13839
rect 41723 13873 41757 13889
rect 41723 13823 41757 13839
rect 1741 13537 1775 13553
rect 1741 13487 1775 13503
rect 41723 13537 41757 13553
rect 41723 13487 41757 13503
rect 1741 13201 1775 13217
rect 1741 13151 1775 13167
rect 41723 13201 41757 13217
rect 41723 13151 41757 13167
rect 1741 12865 1775 12881
rect 1741 12815 1775 12831
rect 41723 12865 41757 12881
rect 41723 12815 41757 12831
rect 1741 12529 1775 12545
rect 1741 12479 1775 12495
rect 41723 12529 41757 12545
rect 41723 12479 41757 12495
rect 1741 12193 1775 12209
rect 1741 12143 1775 12159
rect 41723 12193 41757 12209
rect 41723 12143 41757 12159
rect 1741 11857 1775 11873
rect 1741 11807 1775 11823
rect 41723 11857 41757 11873
rect 41723 11807 41757 11823
rect 1741 11521 1775 11537
rect 1741 11471 1775 11487
rect 41723 11521 41757 11537
rect 41723 11471 41757 11487
rect 1741 11185 1775 11201
rect 1741 11135 1775 11151
rect 41723 11185 41757 11201
rect 41723 11135 41757 11151
rect 1741 10849 1775 10865
rect 1741 10799 1775 10815
rect 41723 10849 41757 10865
rect 41723 10799 41757 10815
rect 1741 10513 1775 10529
rect 1741 10463 1775 10479
rect 41723 10513 41757 10529
rect 41723 10463 41757 10479
rect 1741 10177 1775 10193
rect 1741 10127 1775 10143
rect 41723 10177 41757 10193
rect 41723 10127 41757 10143
rect 1741 9841 1775 9857
rect 1741 9791 1775 9807
rect 41723 9841 41757 9857
rect 41723 9791 41757 9807
rect 1741 9505 1775 9521
rect 1741 9455 1775 9471
rect 41723 9505 41757 9521
rect 41723 9455 41757 9471
rect 1741 9169 1775 9185
rect 1741 9119 1775 9135
rect 41723 9169 41757 9185
rect 41723 9119 41757 9135
rect 1741 8833 1775 8849
rect 1741 8783 1775 8799
rect 41723 8833 41757 8849
rect 41723 8783 41757 8799
rect 1741 8497 1775 8513
rect 1741 8447 1775 8463
rect 41723 8497 41757 8513
rect 41723 8447 41757 8463
rect 1741 8161 1775 8177
rect 1741 8111 1775 8127
rect 41723 8161 41757 8177
rect 41723 8111 41757 8127
rect 1741 7825 1775 7841
rect 1741 7775 1775 7791
rect 41723 7825 41757 7841
rect 41723 7775 41757 7791
rect 1741 7489 1775 7505
rect 1741 7439 1775 7455
rect 41723 7489 41757 7505
rect 41723 7439 41757 7455
rect 1741 7153 1775 7169
rect 1741 7103 1775 7119
rect 41723 7153 41757 7169
rect 41723 7103 41757 7119
rect 1741 6817 1775 6833
rect 1741 6767 1775 6783
rect 41723 6817 41757 6833
rect 41723 6767 41757 6783
rect 1741 6481 1775 6497
rect 1741 6431 1775 6447
rect 41723 6481 41757 6497
rect 41723 6431 41757 6447
rect 1741 6145 1775 6161
rect 1741 6095 1775 6111
rect 41723 6145 41757 6161
rect 41723 6095 41757 6111
rect 1741 5809 1775 5825
rect 1741 5759 1775 5775
rect 41723 5809 41757 5825
rect 41723 5759 41757 5775
rect 1741 5473 1775 5489
rect 1741 5423 1775 5439
rect 41723 5473 41757 5489
rect 41723 5423 41757 5439
rect 1741 5137 1775 5153
rect 1741 5087 1775 5103
rect 41723 5137 41757 5153
rect 41723 5087 41757 5103
rect 1741 4801 1775 4817
rect 1741 4751 1775 4767
rect 41723 4801 41757 4817
rect 41723 4751 41757 4767
rect 1741 4465 1775 4481
rect 1741 4415 1775 4431
rect 41723 4465 41757 4481
rect 41723 4415 41757 4431
rect 1741 4129 1775 4145
rect 1741 4079 1775 4095
rect 41723 4129 41757 4145
rect 41723 4079 41757 4095
rect 1741 3793 1775 3809
rect 1741 3743 1775 3759
rect 41723 3793 41757 3809
rect 41723 3743 41757 3759
rect 1741 3457 1775 3473
rect 1741 3407 1775 3423
rect 41723 3457 41757 3473
rect 41723 3407 41757 3423
rect 1741 3121 1775 3137
rect 1741 3071 1775 3087
rect 41723 3121 41757 3137
rect 41723 3071 41757 3087
rect 1741 2785 1775 2801
rect 1741 2735 1775 2751
rect 41723 2785 41757 2801
rect 41723 2735 41757 2751
rect 1741 2449 1775 2465
rect 1741 2399 1775 2415
rect 41723 2449 41757 2465
rect 41723 2399 41757 2415
rect 1741 2113 1775 2129
rect 1741 2063 1775 2079
rect 41723 2113 41757 2129
rect 41723 2063 41757 2079
rect 2077 1777 2111 1793
rect 2077 1727 2111 1743
rect 2413 1777 2447 1793
rect 2413 1727 2447 1743
rect 2749 1777 2783 1793
rect 2749 1727 2783 1743
rect 3085 1777 3119 1793
rect 3085 1727 3119 1743
rect 3421 1777 3455 1793
rect 3421 1727 3455 1743
rect 3757 1777 3791 1793
rect 3757 1727 3791 1743
rect 4093 1777 4127 1793
rect 4093 1727 4127 1743
rect 4429 1777 4463 1793
rect 4429 1727 4463 1743
rect 4765 1777 4799 1793
rect 4765 1727 4799 1743
rect 5101 1777 5135 1793
rect 5101 1727 5135 1743
rect 5437 1777 5471 1793
rect 5437 1727 5471 1743
rect 5773 1777 5807 1793
rect 5773 1727 5807 1743
rect 6109 1777 6143 1793
rect 6109 1727 6143 1743
rect 6445 1777 6479 1793
rect 6445 1727 6479 1743
rect 6781 1777 6815 1793
rect 6781 1727 6815 1743
rect 7117 1777 7151 1793
rect 7117 1727 7151 1743
rect 7453 1777 7487 1793
rect 7453 1727 7487 1743
rect 7789 1777 7823 1793
rect 7789 1727 7823 1743
rect 8125 1777 8159 1793
rect 8125 1727 8159 1743
rect 8461 1777 8495 1793
rect 8461 1727 8495 1743
rect 8797 1777 8831 1793
rect 8797 1727 8831 1743
rect 9133 1777 9167 1793
rect 9133 1727 9167 1743
rect 9469 1777 9503 1793
rect 9469 1727 9503 1743
rect 9805 1777 9839 1793
rect 9805 1727 9839 1743
rect 10141 1777 10175 1793
rect 10141 1727 10175 1743
rect 10477 1777 10511 1793
rect 10477 1727 10511 1743
rect 10813 1777 10847 1793
rect 10813 1727 10847 1743
rect 11149 1777 11183 1793
rect 11149 1727 11183 1743
rect 11485 1777 11519 1793
rect 11485 1727 11519 1743
rect 11821 1777 11855 1793
rect 11821 1727 11855 1743
rect 12157 1777 12191 1793
rect 12157 1727 12191 1743
rect 12493 1777 12527 1793
rect 12493 1727 12527 1743
rect 12829 1777 12863 1793
rect 12829 1727 12863 1743
rect 13165 1777 13199 1793
rect 13165 1727 13199 1743
rect 13501 1777 13535 1793
rect 13501 1727 13535 1743
rect 13837 1777 13871 1793
rect 13837 1727 13871 1743
rect 14173 1777 14207 1793
rect 14173 1727 14207 1743
rect 14509 1777 14543 1793
rect 14509 1727 14543 1743
rect 14845 1777 14879 1793
rect 14845 1727 14879 1743
rect 15181 1777 15215 1793
rect 15181 1727 15215 1743
rect 15517 1777 15551 1793
rect 15517 1727 15551 1743
rect 15853 1777 15887 1793
rect 15853 1727 15887 1743
rect 16189 1777 16223 1793
rect 16189 1727 16223 1743
rect 16525 1777 16559 1793
rect 16525 1727 16559 1743
rect 16861 1777 16895 1793
rect 16861 1727 16895 1743
rect 17197 1777 17231 1793
rect 17197 1727 17231 1743
rect 17533 1777 17567 1793
rect 17533 1727 17567 1743
rect 17869 1777 17903 1793
rect 17869 1727 17903 1743
rect 18205 1777 18239 1793
rect 18205 1727 18239 1743
rect 18541 1777 18575 1793
rect 18541 1727 18575 1743
rect 18877 1777 18911 1793
rect 18877 1727 18911 1743
rect 19213 1777 19247 1793
rect 19213 1727 19247 1743
rect 19549 1777 19583 1793
rect 19549 1727 19583 1743
rect 19885 1777 19919 1793
rect 19885 1727 19919 1743
rect 20221 1777 20255 1793
rect 20221 1727 20255 1743
rect 20557 1777 20591 1793
rect 20557 1727 20591 1743
rect 20893 1777 20927 1793
rect 20893 1727 20927 1743
rect 21229 1777 21263 1793
rect 21229 1727 21263 1743
rect 21565 1777 21599 1793
rect 21565 1727 21599 1743
rect 21901 1777 21935 1793
rect 21901 1727 21935 1743
rect 22237 1777 22271 1793
rect 22237 1727 22271 1743
rect 22573 1777 22607 1793
rect 22573 1727 22607 1743
rect 22909 1777 22943 1793
rect 22909 1727 22943 1743
rect 23245 1777 23279 1793
rect 23245 1727 23279 1743
rect 23581 1777 23615 1793
rect 23581 1727 23615 1743
rect 23917 1777 23951 1793
rect 23917 1727 23951 1743
rect 24253 1777 24287 1793
rect 24253 1727 24287 1743
rect 24589 1777 24623 1793
rect 24589 1727 24623 1743
rect 24925 1777 24959 1793
rect 24925 1727 24959 1743
rect 25261 1777 25295 1793
rect 25261 1727 25295 1743
rect 25597 1777 25631 1793
rect 25597 1727 25631 1743
rect 25933 1777 25967 1793
rect 25933 1727 25967 1743
rect 26269 1777 26303 1793
rect 26269 1727 26303 1743
rect 26605 1777 26639 1793
rect 26605 1727 26639 1743
rect 26941 1777 26975 1793
rect 26941 1727 26975 1743
rect 27277 1777 27311 1793
rect 27277 1727 27311 1743
rect 27613 1777 27647 1793
rect 27613 1727 27647 1743
rect 27949 1777 27983 1793
rect 27949 1727 27983 1743
rect 28285 1777 28319 1793
rect 28285 1727 28319 1743
rect 28621 1777 28655 1793
rect 28621 1727 28655 1743
rect 28957 1777 28991 1793
rect 28957 1727 28991 1743
rect 29293 1777 29327 1793
rect 29293 1727 29327 1743
rect 29629 1777 29663 1793
rect 29629 1727 29663 1743
rect 29965 1777 29999 1793
rect 29965 1727 29999 1743
rect 30301 1777 30335 1793
rect 30301 1727 30335 1743
rect 30637 1777 30671 1793
rect 30637 1727 30671 1743
rect 30973 1777 31007 1793
rect 30973 1727 31007 1743
rect 31309 1777 31343 1793
rect 31309 1727 31343 1743
rect 31645 1777 31679 1793
rect 31645 1727 31679 1743
rect 31981 1777 32015 1793
rect 31981 1727 32015 1743
rect 32317 1777 32351 1793
rect 32317 1727 32351 1743
rect 32653 1777 32687 1793
rect 32653 1727 32687 1743
rect 32989 1777 33023 1793
rect 32989 1727 33023 1743
rect 33325 1777 33359 1793
rect 33325 1727 33359 1743
rect 33661 1777 33695 1793
rect 33661 1727 33695 1743
rect 33997 1777 34031 1793
rect 33997 1727 34031 1743
rect 34333 1777 34367 1793
rect 34333 1727 34367 1743
rect 34669 1777 34703 1793
rect 34669 1727 34703 1743
rect 35005 1777 35039 1793
rect 35005 1727 35039 1743
rect 35341 1777 35375 1793
rect 35341 1727 35375 1743
rect 35677 1777 35711 1793
rect 35677 1727 35711 1743
rect 36013 1777 36047 1793
rect 36013 1727 36047 1743
rect 36349 1777 36383 1793
rect 36349 1727 36383 1743
rect 36685 1777 36719 1793
rect 36685 1727 36719 1743
rect 37021 1777 37055 1793
rect 37021 1727 37055 1743
rect 37357 1777 37391 1793
rect 37357 1727 37391 1743
rect 37693 1777 37727 1793
rect 37693 1727 37727 1743
rect 38029 1777 38063 1793
rect 38029 1727 38063 1743
rect 38365 1777 38399 1793
rect 38365 1727 38399 1743
rect 38701 1777 38735 1793
rect 38701 1727 38735 1743
rect 39037 1777 39071 1793
rect 39037 1727 39071 1743
rect 39373 1777 39407 1793
rect 39373 1727 39407 1743
rect 39709 1777 39743 1793
rect 39709 1727 39743 1743
rect 40045 1777 40079 1793
rect 40045 1727 40079 1743
rect 40381 1777 40415 1793
rect 40381 1727 40415 1743
rect 40717 1777 40751 1793
rect 40717 1727 40751 1743
rect 41053 1777 41087 1793
rect 41053 1727 41087 1743
<< viali >>
rect 2077 31367 2111 31401
rect 2413 31367 2447 31401
rect 2749 31367 2783 31401
rect 3085 31367 3119 31401
rect 3421 31367 3455 31401
rect 3757 31367 3791 31401
rect 4093 31367 4127 31401
rect 4429 31367 4463 31401
rect 4765 31367 4799 31401
rect 5101 31367 5135 31401
rect 5437 31367 5471 31401
rect 5773 31367 5807 31401
rect 6109 31367 6143 31401
rect 6445 31367 6479 31401
rect 6781 31367 6815 31401
rect 7117 31367 7151 31401
rect 7453 31367 7487 31401
rect 7789 31367 7823 31401
rect 8125 31367 8159 31401
rect 8461 31367 8495 31401
rect 8797 31367 8831 31401
rect 9133 31367 9167 31401
rect 9469 31367 9503 31401
rect 9805 31367 9839 31401
rect 10141 31367 10175 31401
rect 10477 31367 10511 31401
rect 10813 31367 10847 31401
rect 11149 31367 11183 31401
rect 11485 31367 11519 31401
rect 11821 31367 11855 31401
rect 12157 31367 12191 31401
rect 12493 31367 12527 31401
rect 12829 31367 12863 31401
rect 13165 31367 13199 31401
rect 13501 31367 13535 31401
rect 13837 31367 13871 31401
rect 14173 31367 14207 31401
rect 14509 31367 14543 31401
rect 14845 31367 14879 31401
rect 15181 31367 15215 31401
rect 15517 31367 15551 31401
rect 15853 31367 15887 31401
rect 16189 31367 16223 31401
rect 16525 31367 16559 31401
rect 16861 31367 16895 31401
rect 17197 31367 17231 31401
rect 17533 31367 17567 31401
rect 17869 31367 17903 31401
rect 18205 31367 18239 31401
rect 18541 31367 18575 31401
rect 18877 31367 18911 31401
rect 19213 31367 19247 31401
rect 19549 31367 19583 31401
rect 19885 31367 19919 31401
rect 20221 31367 20255 31401
rect 20557 31367 20591 31401
rect 20893 31367 20927 31401
rect 21229 31367 21263 31401
rect 21565 31367 21599 31401
rect 21901 31367 21935 31401
rect 22237 31367 22271 31401
rect 22573 31367 22607 31401
rect 22909 31367 22943 31401
rect 23245 31367 23279 31401
rect 23581 31367 23615 31401
rect 23917 31367 23951 31401
rect 24253 31367 24287 31401
rect 24589 31367 24623 31401
rect 24925 31367 24959 31401
rect 25261 31367 25295 31401
rect 25597 31367 25631 31401
rect 25933 31367 25967 31401
rect 26269 31367 26303 31401
rect 26605 31367 26639 31401
rect 26941 31367 26975 31401
rect 27277 31367 27311 31401
rect 27613 31367 27647 31401
rect 27949 31367 27983 31401
rect 28285 31367 28319 31401
rect 28621 31367 28655 31401
rect 28957 31367 28991 31401
rect 29293 31367 29327 31401
rect 29629 31367 29663 31401
rect 29965 31367 29999 31401
rect 30301 31367 30335 31401
rect 30637 31367 30671 31401
rect 30973 31367 31007 31401
rect 31309 31367 31343 31401
rect 31645 31367 31679 31401
rect 31981 31367 32015 31401
rect 32317 31367 32351 31401
rect 32653 31367 32687 31401
rect 32989 31367 33023 31401
rect 33325 31367 33359 31401
rect 33661 31367 33695 31401
rect 33997 31367 34031 31401
rect 34333 31367 34367 31401
rect 34669 31367 34703 31401
rect 35005 31367 35039 31401
rect 35341 31367 35375 31401
rect 35677 31367 35711 31401
rect 36013 31367 36047 31401
rect 36349 31367 36383 31401
rect 36685 31367 36719 31401
rect 37021 31367 37055 31401
rect 37357 31367 37391 31401
rect 37693 31367 37727 31401
rect 38029 31367 38063 31401
rect 38365 31367 38399 31401
rect 38701 31367 38735 31401
rect 39037 31367 39071 31401
rect 39373 31367 39407 31401
rect 39709 31367 39743 31401
rect 40045 31367 40079 31401
rect 40381 31367 40415 31401
rect 40717 31367 40751 31401
rect 41053 31367 41087 31401
rect 1741 30975 1775 31009
rect 41723 30975 41757 31009
rect 1741 30639 1775 30673
rect 41723 30639 41757 30673
rect 1741 30303 1775 30337
rect 41723 30303 41757 30337
rect 1741 29967 1775 30001
rect 41723 29967 41757 30001
rect 1741 29631 1775 29665
rect 41723 29631 41757 29665
rect 1741 29295 1775 29329
rect 41723 29295 41757 29329
rect 1741 28959 1775 28993
rect 41723 28959 41757 28993
rect 1741 28623 1775 28657
rect 41723 28623 41757 28657
rect 1741 28287 1775 28321
rect 41723 28287 41757 28321
rect 1741 27951 1775 27985
rect 41723 27951 41757 27985
rect 1741 27615 1775 27649
rect 41723 27615 41757 27649
rect 1741 27279 1775 27313
rect 41723 27279 41757 27313
rect 1741 26943 1775 26977
rect 41723 26943 41757 26977
rect 1741 26607 1775 26641
rect 41723 26607 41757 26641
rect 1741 26271 1775 26305
rect 41723 26271 41757 26305
rect 1741 25935 1775 25969
rect 41723 25935 41757 25969
rect 1741 25599 1775 25633
rect 41723 25599 41757 25633
rect 1741 25263 1775 25297
rect 41723 25263 41757 25297
rect 1741 24927 1775 24961
rect 41723 24927 41757 24961
rect 1741 24591 1775 24625
rect 41723 24591 41757 24625
rect 1741 24255 1775 24289
rect 41723 24255 41757 24289
rect 1741 23919 1775 23953
rect 41723 23919 41757 23953
rect 1741 23583 1775 23617
rect 41723 23583 41757 23617
rect 1741 23247 1775 23281
rect 41723 23247 41757 23281
rect 1741 22911 1775 22945
rect 41723 22911 41757 22945
rect 1741 22575 1775 22609
rect 41723 22575 41757 22609
rect 1741 22239 1775 22273
rect 41723 22239 41757 22273
rect 1741 21903 1775 21937
rect 41723 21903 41757 21937
rect 1741 21567 1775 21601
rect 41723 21567 41757 21601
rect 1741 21231 1775 21265
rect 41723 21231 41757 21265
rect 1741 20895 1775 20929
rect 41723 20895 41757 20929
rect 1741 20559 1775 20593
rect 41723 20559 41757 20593
rect 1741 20223 1775 20257
rect 41723 20223 41757 20257
rect 1741 19887 1775 19921
rect 41723 19887 41757 19921
rect 1741 19551 1775 19585
rect 41723 19551 41757 19585
rect 1741 19215 1775 19249
rect 41723 19215 41757 19249
rect 1741 18879 1775 18913
rect 41723 18879 41757 18913
rect 1741 18543 1775 18577
rect 41723 18543 41757 18577
rect 1741 18207 1775 18241
rect 41723 18207 41757 18241
rect 1741 17871 1775 17905
rect 41723 17871 41757 17905
rect 1741 17535 1775 17569
rect 41723 17535 41757 17569
rect 1741 17199 1775 17233
rect 41723 17199 41757 17233
rect 1741 16863 1775 16897
rect 41723 16863 41757 16897
rect 1741 16527 1775 16561
rect 41723 16527 41757 16561
rect 1741 16191 1775 16225
rect 41723 16191 41757 16225
rect 1741 15855 1775 15889
rect 41723 15855 41757 15889
rect 1741 15519 1775 15553
rect 41723 15519 41757 15553
rect 1741 15183 1775 15217
rect 41723 15183 41757 15217
rect 1741 14847 1775 14881
rect 41723 14847 41757 14881
rect 1741 14511 1775 14545
rect 41723 14511 41757 14545
rect 1741 14175 1775 14209
rect 41723 14175 41757 14209
rect 1741 13839 1775 13873
rect 41723 13839 41757 13873
rect 1741 13503 1775 13537
rect 41723 13503 41757 13537
rect 1741 13167 1775 13201
rect 41723 13167 41757 13201
rect 1741 12831 1775 12865
rect 41723 12831 41757 12865
rect 1741 12495 1775 12529
rect 41723 12495 41757 12529
rect 1741 12159 1775 12193
rect 41723 12159 41757 12193
rect 1741 11823 1775 11857
rect 41723 11823 41757 11857
rect 1741 11487 1775 11521
rect 41723 11487 41757 11521
rect 1741 11151 1775 11185
rect 41723 11151 41757 11185
rect 1741 10815 1775 10849
rect 41723 10815 41757 10849
rect 1741 10479 1775 10513
rect 41723 10479 41757 10513
rect 1741 10143 1775 10177
rect 41723 10143 41757 10177
rect 1741 9807 1775 9841
rect 41723 9807 41757 9841
rect 1741 9471 1775 9505
rect 41723 9471 41757 9505
rect 1741 9135 1775 9169
rect 41723 9135 41757 9169
rect 1741 8799 1775 8833
rect 41723 8799 41757 8833
rect 1741 8463 1775 8497
rect 41723 8463 41757 8497
rect 1741 8127 1775 8161
rect 41723 8127 41757 8161
rect 1741 7791 1775 7825
rect 41723 7791 41757 7825
rect 1741 7455 1775 7489
rect 41723 7455 41757 7489
rect 1741 7119 1775 7153
rect 41723 7119 41757 7153
rect 1741 6783 1775 6817
rect 41723 6783 41757 6817
rect 1741 6447 1775 6481
rect 41723 6447 41757 6481
rect 1741 6111 1775 6145
rect 41723 6111 41757 6145
rect 1741 5775 1775 5809
rect 41723 5775 41757 5809
rect 1741 5439 1775 5473
rect 41723 5439 41757 5473
rect 1741 5103 1775 5137
rect 41723 5103 41757 5137
rect 1741 4767 1775 4801
rect 41723 4767 41757 4801
rect 1741 4431 1775 4465
rect 41723 4431 41757 4465
rect 1741 4095 1775 4129
rect 41723 4095 41757 4129
rect 1741 3759 1775 3793
rect 41723 3759 41757 3793
rect 1741 3423 1775 3457
rect 41723 3423 41757 3457
rect 1741 3087 1775 3121
rect 41723 3087 41757 3121
rect 1741 2751 1775 2785
rect 41723 2751 41757 2785
rect 1741 2415 1775 2449
rect 41723 2415 41757 2449
rect 1741 2079 1775 2113
rect 41723 2079 41757 2113
rect 2077 1743 2111 1777
rect 2413 1743 2447 1777
rect 2749 1743 2783 1777
rect 3085 1743 3119 1777
rect 3421 1743 3455 1777
rect 3757 1743 3791 1777
rect 4093 1743 4127 1777
rect 4429 1743 4463 1777
rect 4765 1743 4799 1777
rect 5101 1743 5135 1777
rect 5437 1743 5471 1777
rect 5773 1743 5807 1777
rect 6109 1743 6143 1777
rect 6445 1743 6479 1777
rect 6781 1743 6815 1777
rect 7117 1743 7151 1777
rect 7453 1743 7487 1777
rect 7789 1743 7823 1777
rect 8125 1743 8159 1777
rect 8461 1743 8495 1777
rect 8797 1743 8831 1777
rect 9133 1743 9167 1777
rect 9469 1743 9503 1777
rect 9805 1743 9839 1777
rect 10141 1743 10175 1777
rect 10477 1743 10511 1777
rect 10813 1743 10847 1777
rect 11149 1743 11183 1777
rect 11485 1743 11519 1777
rect 11821 1743 11855 1777
rect 12157 1743 12191 1777
rect 12493 1743 12527 1777
rect 12829 1743 12863 1777
rect 13165 1743 13199 1777
rect 13501 1743 13535 1777
rect 13837 1743 13871 1777
rect 14173 1743 14207 1777
rect 14509 1743 14543 1777
rect 14845 1743 14879 1777
rect 15181 1743 15215 1777
rect 15517 1743 15551 1777
rect 15853 1743 15887 1777
rect 16189 1743 16223 1777
rect 16525 1743 16559 1777
rect 16861 1743 16895 1777
rect 17197 1743 17231 1777
rect 17533 1743 17567 1777
rect 17869 1743 17903 1777
rect 18205 1743 18239 1777
rect 18541 1743 18575 1777
rect 18877 1743 18911 1777
rect 19213 1743 19247 1777
rect 19549 1743 19583 1777
rect 19885 1743 19919 1777
rect 20221 1743 20255 1777
rect 20557 1743 20591 1777
rect 20893 1743 20927 1777
rect 21229 1743 21263 1777
rect 21565 1743 21599 1777
rect 21901 1743 21935 1777
rect 22237 1743 22271 1777
rect 22573 1743 22607 1777
rect 22909 1743 22943 1777
rect 23245 1743 23279 1777
rect 23581 1743 23615 1777
rect 23917 1743 23951 1777
rect 24253 1743 24287 1777
rect 24589 1743 24623 1777
rect 24925 1743 24959 1777
rect 25261 1743 25295 1777
rect 25597 1743 25631 1777
rect 25933 1743 25967 1777
rect 26269 1743 26303 1777
rect 26605 1743 26639 1777
rect 26941 1743 26975 1777
rect 27277 1743 27311 1777
rect 27613 1743 27647 1777
rect 27949 1743 27983 1777
rect 28285 1743 28319 1777
rect 28621 1743 28655 1777
rect 28957 1743 28991 1777
rect 29293 1743 29327 1777
rect 29629 1743 29663 1777
rect 29965 1743 29999 1777
rect 30301 1743 30335 1777
rect 30637 1743 30671 1777
rect 30973 1743 31007 1777
rect 31309 1743 31343 1777
rect 31645 1743 31679 1777
rect 31981 1743 32015 1777
rect 32317 1743 32351 1777
rect 32653 1743 32687 1777
rect 32989 1743 33023 1777
rect 33325 1743 33359 1777
rect 33661 1743 33695 1777
rect 33997 1743 34031 1777
rect 34333 1743 34367 1777
rect 34669 1743 34703 1777
rect 35005 1743 35039 1777
rect 35341 1743 35375 1777
rect 35677 1743 35711 1777
rect 36013 1743 36047 1777
rect 36349 1743 36383 1777
rect 36685 1743 36719 1777
rect 37021 1743 37055 1777
rect 37357 1743 37391 1777
rect 37693 1743 37727 1777
rect 38029 1743 38063 1777
rect 38365 1743 38399 1777
rect 38701 1743 38735 1777
rect 39037 1743 39071 1777
rect 39373 1743 39407 1777
rect 39709 1743 39743 1777
rect 40045 1743 40079 1777
rect 40381 1743 40415 1777
rect 40717 1743 40751 1777
rect 41053 1743 41087 1777
<< metal1 >>
rect 1646 31410 41852 31496
rect 1646 31358 2068 31410
rect 2120 31401 3748 31410
rect 3800 31401 5428 31410
rect 5480 31401 7108 31410
rect 7160 31401 8788 31410
rect 8840 31401 10468 31410
rect 10520 31401 12148 31410
rect 12200 31401 13828 31410
rect 13880 31401 15508 31410
rect 15560 31401 17188 31410
rect 17240 31401 18868 31410
rect 18920 31401 20548 31410
rect 20600 31401 22228 31410
rect 22280 31401 23908 31410
rect 23960 31401 25588 31410
rect 25640 31401 27268 31410
rect 27320 31401 28948 31410
rect 29000 31401 30628 31410
rect 30680 31401 32308 31410
rect 32360 31401 33988 31410
rect 34040 31401 35668 31410
rect 35720 31401 37348 31410
rect 37400 31401 39028 31410
rect 39080 31401 40708 31410
rect 40760 31401 41852 31410
rect 2120 31367 2413 31401
rect 2447 31367 2749 31401
rect 2783 31367 3085 31401
rect 3119 31367 3421 31401
rect 3455 31367 3748 31401
rect 3800 31367 4093 31401
rect 4127 31367 4429 31401
rect 4463 31367 4765 31401
rect 4799 31367 5101 31401
rect 5135 31367 5428 31401
rect 5480 31367 5773 31401
rect 5807 31367 6109 31401
rect 6143 31367 6445 31401
rect 6479 31367 6781 31401
rect 6815 31367 7108 31401
rect 7160 31367 7453 31401
rect 7487 31367 7789 31401
rect 7823 31367 8125 31401
rect 8159 31367 8461 31401
rect 8495 31367 8788 31401
rect 8840 31367 9133 31401
rect 9167 31367 9469 31401
rect 9503 31367 9805 31401
rect 9839 31367 10141 31401
rect 10175 31367 10468 31401
rect 10520 31367 10813 31401
rect 10847 31367 11149 31401
rect 11183 31367 11485 31401
rect 11519 31367 11821 31401
rect 11855 31367 12148 31401
rect 12200 31367 12493 31401
rect 12527 31367 12829 31401
rect 12863 31367 13165 31401
rect 13199 31367 13501 31401
rect 13535 31367 13828 31401
rect 13880 31367 14173 31401
rect 14207 31367 14509 31401
rect 14543 31367 14845 31401
rect 14879 31367 15181 31401
rect 15215 31367 15508 31401
rect 15560 31367 15853 31401
rect 15887 31367 16189 31401
rect 16223 31367 16525 31401
rect 16559 31367 16861 31401
rect 16895 31367 17188 31401
rect 17240 31367 17533 31401
rect 17567 31367 17869 31401
rect 17903 31367 18205 31401
rect 18239 31367 18541 31401
rect 18575 31367 18868 31401
rect 18920 31367 19213 31401
rect 19247 31367 19549 31401
rect 19583 31367 19885 31401
rect 19919 31367 20221 31401
rect 20255 31367 20548 31401
rect 20600 31367 20893 31401
rect 20927 31367 21229 31401
rect 21263 31367 21565 31401
rect 21599 31367 21901 31401
rect 21935 31367 22228 31401
rect 22280 31367 22573 31401
rect 22607 31367 22909 31401
rect 22943 31367 23245 31401
rect 23279 31367 23581 31401
rect 23615 31367 23908 31401
rect 23960 31367 24253 31401
rect 24287 31367 24589 31401
rect 24623 31367 24925 31401
rect 24959 31367 25261 31401
rect 25295 31367 25588 31401
rect 25640 31367 25933 31401
rect 25967 31367 26269 31401
rect 26303 31367 26605 31401
rect 26639 31367 26941 31401
rect 26975 31367 27268 31401
rect 27320 31367 27613 31401
rect 27647 31367 27949 31401
rect 27983 31367 28285 31401
rect 28319 31367 28621 31401
rect 28655 31367 28948 31401
rect 29000 31367 29293 31401
rect 29327 31367 29629 31401
rect 29663 31367 29965 31401
rect 29999 31367 30301 31401
rect 30335 31367 30628 31401
rect 30680 31367 30973 31401
rect 31007 31367 31309 31401
rect 31343 31367 31645 31401
rect 31679 31367 31981 31401
rect 32015 31367 32308 31401
rect 32360 31367 32653 31401
rect 32687 31367 32989 31401
rect 33023 31367 33325 31401
rect 33359 31367 33661 31401
rect 33695 31367 33988 31401
rect 34040 31367 34333 31401
rect 34367 31367 34669 31401
rect 34703 31367 35005 31401
rect 35039 31367 35341 31401
rect 35375 31367 35668 31401
rect 35720 31367 36013 31401
rect 36047 31367 36349 31401
rect 36383 31367 36685 31401
rect 36719 31367 37021 31401
rect 37055 31367 37348 31401
rect 37400 31367 37693 31401
rect 37727 31367 38029 31401
rect 38063 31367 38365 31401
rect 38399 31367 38701 31401
rect 38735 31367 39028 31401
rect 39080 31367 39373 31401
rect 39407 31367 39709 31401
rect 39743 31367 40045 31401
rect 40079 31367 40381 31401
rect 40415 31367 40708 31401
rect 40760 31367 41053 31401
rect 41087 31367 41852 31401
rect 2120 31358 3748 31367
rect 3800 31358 5428 31367
rect 5480 31358 7108 31367
rect 7160 31358 8788 31367
rect 8840 31358 10468 31367
rect 10520 31358 12148 31367
rect 12200 31358 13828 31367
rect 13880 31358 15508 31367
rect 15560 31358 17188 31367
rect 17240 31358 18868 31367
rect 18920 31358 20548 31367
rect 20600 31358 22228 31367
rect 22280 31358 23908 31367
rect 23960 31358 25588 31367
rect 25640 31358 27268 31367
rect 27320 31358 28948 31367
rect 29000 31358 30628 31367
rect 30680 31358 32308 31367
rect 32360 31358 33988 31367
rect 34040 31358 35668 31367
rect 35720 31358 37348 31367
rect 37400 31358 39028 31367
rect 39080 31358 40708 31367
rect 40760 31358 41852 31367
rect 1646 31272 41852 31358
rect 1726 30966 1732 31018
rect 1784 30966 1790 31018
rect 41708 30966 41714 31018
rect 41766 30966 41772 31018
rect 1726 30630 1732 30682
rect 1784 30630 1790 30682
rect 41708 30630 41714 30682
rect 41766 30630 41772 30682
rect 1726 30294 1732 30346
rect 1784 30294 1790 30346
rect 41708 30294 41714 30346
rect 41766 30294 41772 30346
rect 1726 29958 1732 30010
rect 1784 29958 1790 30010
rect 41708 29958 41714 30010
rect 41766 29958 41772 30010
rect 1726 29622 1732 29674
rect 1784 29622 1790 29674
rect 41708 29622 41714 29674
rect 41766 29622 41772 29674
rect 1726 29286 1732 29338
rect 1784 29286 1790 29338
rect 41708 29286 41714 29338
rect 41766 29286 41772 29338
rect 1726 28950 1732 29002
rect 1784 28950 1790 29002
rect 41708 28950 41714 29002
rect 41766 28950 41772 29002
rect 1726 28614 1732 28666
rect 1784 28614 1790 28666
rect 41708 28614 41714 28666
rect 41766 28614 41772 28666
rect 1726 28278 1732 28330
rect 1784 28278 1790 28330
rect 41708 28278 41714 28330
rect 41766 28278 41772 28330
rect 1726 27942 1732 27994
rect 1784 27942 1790 27994
rect 41708 27942 41714 27994
rect 41766 27942 41772 27994
rect 1726 27606 1732 27658
rect 1784 27606 1790 27658
rect 41708 27606 41714 27658
rect 41766 27606 41772 27658
rect 1726 27270 1732 27322
rect 1784 27270 1790 27322
rect 41708 27270 41714 27322
rect 41766 27270 41772 27322
rect 1726 26934 1732 26986
rect 1784 26934 1790 26986
rect 41708 26934 41714 26986
rect 41766 26934 41772 26986
rect 1726 26598 1732 26650
rect 1784 26598 1790 26650
rect 41708 26598 41714 26650
rect 41766 26598 41772 26650
rect 1726 26262 1732 26314
rect 1784 26262 1790 26314
rect 41708 26262 41714 26314
rect 41766 26262 41772 26314
rect 9935 26137 9941 26189
rect 9993 26137 9999 26189
rect 1726 25926 1732 25978
rect 1784 25926 1790 25978
rect 1726 25590 1732 25642
rect 1784 25590 1790 25642
rect 1726 25254 1732 25306
rect 1784 25254 1790 25306
rect 1726 24918 1732 24970
rect 1784 24918 1790 24970
rect 1726 24582 1732 24634
rect 1784 24582 1790 24634
rect 9855 24579 9861 24631
rect 9913 24579 9919 24631
rect 1726 24246 1732 24298
rect 1784 24246 1790 24298
rect 1726 23910 1732 23962
rect 1784 23910 1790 23962
rect 1726 23574 1732 23626
rect 1784 23574 1790 23626
rect 9775 23309 9781 23361
rect 9833 23309 9839 23361
rect 1726 23238 1732 23290
rect 1784 23238 1790 23290
rect 1726 22902 1732 22954
rect 1784 22902 1790 22954
rect 1726 22566 1732 22618
rect 1784 22566 1790 22618
rect 1726 22230 1732 22282
rect 1784 22230 1790 22282
rect 1726 21894 1732 21946
rect 1784 21894 1790 21946
rect 9695 21751 9701 21803
rect 9753 21751 9759 21803
rect 1726 21558 1732 21610
rect 1784 21558 1790 21610
rect 1726 21222 1732 21274
rect 1784 21222 1790 21274
rect 1726 20886 1732 20938
rect 1784 20886 1790 20938
rect 1726 20550 1732 20602
rect 1784 20550 1790 20602
rect 1726 20214 1732 20266
rect 1784 20214 1790 20266
rect 1726 19878 1732 19930
rect 1784 19878 1790 19930
rect 1726 19542 1732 19594
rect 1784 19542 1790 19594
rect 1726 19206 1732 19258
rect 1784 19206 1790 19258
rect 1726 18870 1732 18922
rect 1784 18870 1790 18922
rect 1726 18534 1732 18586
rect 1784 18534 1790 18586
rect 1726 18198 1732 18250
rect 1784 18198 1790 18250
rect 1726 17862 1732 17914
rect 1784 17862 1790 17914
rect 1726 17526 1732 17578
rect 1784 17526 1790 17578
rect 1726 17190 1732 17242
rect 1784 17190 1790 17242
rect 1726 16854 1732 16906
rect 1784 16854 1790 16906
rect 9713 16801 9741 21751
rect 9793 16801 9821 23309
rect 9873 16801 9901 24579
rect 9953 16801 9981 26137
rect 41708 25926 41714 25978
rect 41766 25926 41772 25978
rect 41708 25590 41714 25642
rect 41766 25590 41772 25642
rect 19402 25297 19408 25349
rect 19460 25297 19466 25349
rect 20396 25297 20402 25349
rect 20454 25297 20460 25349
rect 20650 25297 20656 25349
rect 20708 25297 20714 25349
rect 21644 25297 21650 25349
rect 21702 25297 21708 25349
rect 21898 25297 21904 25349
rect 21956 25297 21962 25349
rect 22892 25297 22898 25349
rect 22950 25297 22956 25349
rect 23146 25297 23152 25349
rect 23204 25297 23210 25349
rect 24140 25297 24146 25349
rect 24198 25297 24204 25349
rect 41708 25254 41714 25306
rect 41766 25254 41772 25306
rect 41708 24918 41714 24970
rect 41766 24918 41772 24970
rect 41708 24582 41714 24634
rect 41766 24582 41772 24634
rect 41708 24246 41714 24298
rect 41766 24246 41772 24298
rect 41708 23910 41714 23962
rect 41766 23910 41772 23962
rect 41708 23574 41714 23626
rect 41766 23574 41772 23626
rect 41708 23238 41714 23290
rect 41766 23238 41772 23290
rect 41708 22902 41714 22954
rect 41766 22902 41772 22954
rect 41708 22566 41714 22618
rect 41766 22566 41772 22618
rect 41708 22230 41714 22282
rect 41766 22230 41772 22282
rect 41708 21894 41714 21946
rect 41766 21894 41772 21946
rect 41708 21558 41714 21610
rect 41766 21558 41772 21610
rect 41708 21222 41714 21274
rect 41766 21222 41772 21274
rect 41708 20886 41714 20938
rect 41766 20886 41772 20938
rect 41708 20550 41714 20602
rect 41766 20550 41772 20602
rect 41708 20214 41714 20266
rect 41766 20214 41772 20266
rect 41708 19878 41714 19930
rect 41766 19878 41772 19930
rect 41708 19542 41714 19594
rect 41766 19542 41772 19594
rect 41708 19206 41714 19258
rect 41766 19206 41772 19258
rect 41708 18870 41714 18922
rect 41766 18870 41772 18922
rect 41708 18534 41714 18586
rect 41766 18534 41772 18586
rect 41708 18198 41714 18250
rect 41766 18198 41772 18250
rect 41708 17862 41714 17914
rect 41766 17862 41772 17914
rect 41708 17526 41714 17578
rect 41766 17526 41772 17578
rect 41708 17190 41714 17242
rect 41766 17190 41772 17242
rect 41708 16854 41714 16906
rect 41766 16854 41772 16906
rect 1726 16518 1732 16570
rect 1784 16518 1790 16570
rect 1726 16182 1732 16234
rect 1784 16182 1790 16234
rect 1726 15846 1732 15898
rect 1784 15846 1790 15898
rect 1726 15510 1732 15562
rect 1784 15510 1790 15562
rect 1726 15174 1732 15226
rect 1784 15174 1790 15226
rect 1726 14838 1732 14890
rect 1784 14838 1790 14890
rect 1726 14502 1732 14554
rect 1784 14502 1790 14554
rect 1726 14166 1732 14218
rect 1784 14166 1790 14218
rect 1726 13830 1732 13882
rect 1784 13830 1790 13882
rect 1726 13494 1732 13546
rect 1784 13494 1790 13546
rect 1726 13158 1732 13210
rect 1784 13158 1790 13210
rect 1726 12822 1732 12874
rect 1784 12822 1790 12874
rect 1726 12486 1732 12538
rect 1784 12486 1790 12538
rect 1726 12150 1732 12202
rect 1784 12150 1790 12202
rect 1726 11814 1732 11866
rect 1784 11814 1790 11866
rect 1726 11478 1732 11530
rect 1784 11478 1790 11530
rect 1726 11142 1732 11194
rect 1784 11142 1790 11194
rect 1726 10806 1732 10858
rect 1784 10806 1790 10858
rect 19402 10623 19408 10675
rect 19460 10623 19466 10675
rect 20396 10623 20402 10675
rect 20454 10623 20460 10675
rect 20650 10623 20656 10675
rect 20708 10623 20714 10675
rect 21644 10623 21650 10675
rect 21702 10623 21708 10675
rect 21898 10623 21904 10675
rect 21956 10623 21962 10675
rect 22892 10623 22898 10675
rect 22950 10623 22956 10675
rect 23146 10623 23152 10675
rect 23204 10623 23210 10675
rect 24140 10623 24146 10675
rect 24198 10623 24204 10675
rect 1726 10470 1732 10522
rect 1784 10470 1790 10522
rect 1726 10134 1732 10186
rect 1784 10134 1790 10186
rect 1726 9798 1732 9850
rect 1784 9798 1790 9850
rect 33625 9831 33653 16801
rect 33705 11389 33733 16801
rect 33785 12659 33813 16801
rect 33865 14217 33893 16801
rect 41708 16518 41714 16570
rect 41766 16518 41772 16570
rect 41708 16182 41714 16234
rect 41766 16182 41772 16234
rect 41708 15846 41714 15898
rect 41766 15846 41772 15898
rect 41708 15510 41714 15562
rect 41766 15510 41772 15562
rect 41708 15174 41714 15226
rect 41766 15174 41772 15226
rect 41708 14838 41714 14890
rect 41766 14838 41772 14890
rect 41708 14502 41714 14554
rect 41766 14502 41772 14554
rect 33847 14165 33853 14217
rect 33905 14165 33911 14217
rect 41708 14166 41714 14218
rect 41766 14166 41772 14218
rect 41708 13830 41714 13882
rect 41766 13830 41772 13882
rect 41708 13494 41714 13546
rect 41766 13494 41772 13546
rect 41708 13158 41714 13210
rect 41766 13158 41772 13210
rect 41708 12822 41714 12874
rect 41766 12822 41772 12874
rect 33767 12607 33773 12659
rect 33825 12607 33831 12659
rect 41708 12486 41714 12538
rect 41766 12486 41772 12538
rect 41708 12150 41714 12202
rect 41766 12150 41772 12202
rect 41708 11814 41714 11866
rect 41766 11814 41772 11866
rect 41708 11478 41714 11530
rect 41766 11478 41772 11530
rect 33687 11337 33693 11389
rect 33745 11337 33751 11389
rect 41708 11142 41714 11194
rect 41766 11142 41772 11194
rect 41708 10806 41714 10858
rect 41766 10806 41772 10858
rect 41708 10470 41714 10522
rect 41766 10470 41772 10522
rect 41708 10134 41714 10186
rect 41766 10134 41772 10186
rect 33607 9779 33613 9831
rect 33665 9779 33671 9831
rect 41708 9798 41714 9850
rect 41766 9798 41772 9850
rect 1726 9462 1732 9514
rect 1784 9462 1790 9514
rect 41708 9462 41714 9514
rect 41766 9462 41772 9514
rect 1726 9126 1732 9178
rect 1784 9126 1790 9178
rect 41708 9126 41714 9178
rect 41766 9126 41772 9178
rect 1726 8790 1732 8842
rect 1784 8790 1790 8842
rect 41708 8790 41714 8842
rect 41766 8790 41772 8842
rect 1726 8454 1732 8506
rect 1784 8454 1790 8506
rect 41708 8454 41714 8506
rect 41766 8454 41772 8506
rect 1726 8118 1732 8170
rect 1784 8118 1790 8170
rect 41708 8118 41714 8170
rect 41766 8118 41772 8170
rect 1726 7782 1732 7834
rect 1784 7782 1790 7834
rect 41708 7782 41714 7834
rect 41766 7782 41772 7834
rect 1726 7446 1732 7498
rect 1784 7446 1790 7498
rect 41708 7446 41714 7498
rect 41766 7446 41772 7498
rect 1726 7110 1732 7162
rect 1784 7110 1790 7162
rect 41708 7110 41714 7162
rect 41766 7110 41772 7162
rect 1726 6774 1732 6826
rect 1784 6774 1790 6826
rect 41708 6774 41714 6826
rect 41766 6774 41772 6826
rect 1726 6438 1732 6490
rect 1784 6438 1790 6490
rect 41708 6438 41714 6490
rect 41766 6438 41772 6490
rect 1726 6102 1732 6154
rect 1784 6102 1790 6154
rect 41708 6102 41714 6154
rect 41766 6102 41772 6154
rect 1726 5766 1732 5818
rect 1784 5766 1790 5818
rect 41708 5766 41714 5818
rect 41766 5766 41772 5818
rect 1726 5430 1732 5482
rect 1784 5430 1790 5482
rect 41708 5430 41714 5482
rect 41766 5430 41772 5482
rect 1726 5094 1732 5146
rect 1784 5094 1790 5146
rect 41708 5094 41714 5146
rect 41766 5094 41772 5146
rect 1726 4758 1732 4810
rect 1784 4758 1790 4810
rect 41708 4758 41714 4810
rect 41766 4758 41772 4810
rect 1726 4422 1732 4474
rect 1784 4422 1790 4474
rect 41708 4422 41714 4474
rect 41766 4422 41772 4474
rect 1726 4086 1732 4138
rect 1784 4086 1790 4138
rect 41708 4086 41714 4138
rect 41766 4086 41772 4138
rect 1726 3750 1732 3802
rect 1784 3750 1790 3802
rect 41708 3750 41714 3802
rect 41766 3750 41772 3802
rect 1726 3414 1732 3466
rect 1784 3414 1790 3466
rect 41708 3414 41714 3466
rect 41766 3414 41772 3466
rect 1726 3078 1732 3130
rect 1784 3078 1790 3130
rect 41708 3078 41714 3130
rect 41766 3078 41772 3130
rect 1726 2742 1732 2794
rect 1784 2742 1790 2794
rect 41708 2742 41714 2794
rect 41766 2742 41772 2794
rect 1726 2406 1732 2458
rect 1784 2406 1790 2458
rect 41708 2406 41714 2458
rect 41766 2406 41772 2458
rect 1726 2070 1732 2122
rect 1784 2070 1790 2122
rect 41708 2070 41714 2122
rect 41766 2070 41772 2122
rect 1646 1786 41852 1872
rect 1646 1734 2068 1786
rect 2120 1777 3748 1786
rect 3800 1777 5428 1786
rect 5480 1777 7108 1786
rect 7160 1777 8788 1786
rect 8840 1777 10468 1786
rect 10520 1777 12148 1786
rect 12200 1777 13828 1786
rect 13880 1777 15508 1786
rect 15560 1777 17188 1786
rect 17240 1777 18868 1786
rect 18920 1777 20548 1786
rect 20600 1777 22228 1786
rect 22280 1777 23908 1786
rect 23960 1777 25588 1786
rect 25640 1777 27268 1786
rect 27320 1777 28948 1786
rect 29000 1777 30628 1786
rect 30680 1777 32308 1786
rect 32360 1777 33988 1786
rect 34040 1777 35668 1786
rect 35720 1777 37348 1786
rect 37400 1777 39028 1786
rect 39080 1777 40708 1786
rect 40760 1777 41852 1786
rect 2120 1743 2413 1777
rect 2447 1743 2749 1777
rect 2783 1743 3085 1777
rect 3119 1743 3421 1777
rect 3455 1743 3748 1777
rect 3800 1743 4093 1777
rect 4127 1743 4429 1777
rect 4463 1743 4765 1777
rect 4799 1743 5101 1777
rect 5135 1743 5428 1777
rect 5480 1743 5773 1777
rect 5807 1743 6109 1777
rect 6143 1743 6445 1777
rect 6479 1743 6781 1777
rect 6815 1743 7108 1777
rect 7160 1743 7453 1777
rect 7487 1743 7789 1777
rect 7823 1743 8125 1777
rect 8159 1743 8461 1777
rect 8495 1743 8788 1777
rect 8840 1743 9133 1777
rect 9167 1743 9469 1777
rect 9503 1743 9805 1777
rect 9839 1743 10141 1777
rect 10175 1743 10468 1777
rect 10520 1743 10813 1777
rect 10847 1743 11149 1777
rect 11183 1743 11485 1777
rect 11519 1743 11821 1777
rect 11855 1743 12148 1777
rect 12200 1743 12493 1777
rect 12527 1743 12829 1777
rect 12863 1743 13165 1777
rect 13199 1743 13501 1777
rect 13535 1743 13828 1777
rect 13880 1743 14173 1777
rect 14207 1743 14509 1777
rect 14543 1743 14845 1777
rect 14879 1743 15181 1777
rect 15215 1743 15508 1777
rect 15560 1743 15853 1777
rect 15887 1743 16189 1777
rect 16223 1743 16525 1777
rect 16559 1743 16861 1777
rect 16895 1743 17188 1777
rect 17240 1743 17533 1777
rect 17567 1743 17869 1777
rect 17903 1743 18205 1777
rect 18239 1743 18541 1777
rect 18575 1743 18868 1777
rect 18920 1743 19213 1777
rect 19247 1743 19549 1777
rect 19583 1743 19885 1777
rect 19919 1743 20221 1777
rect 20255 1743 20548 1777
rect 20600 1743 20893 1777
rect 20927 1743 21229 1777
rect 21263 1743 21565 1777
rect 21599 1743 21901 1777
rect 21935 1743 22228 1777
rect 22280 1743 22573 1777
rect 22607 1743 22909 1777
rect 22943 1743 23245 1777
rect 23279 1743 23581 1777
rect 23615 1743 23908 1777
rect 23960 1743 24253 1777
rect 24287 1743 24589 1777
rect 24623 1743 24925 1777
rect 24959 1743 25261 1777
rect 25295 1743 25588 1777
rect 25640 1743 25933 1777
rect 25967 1743 26269 1777
rect 26303 1743 26605 1777
rect 26639 1743 26941 1777
rect 26975 1743 27268 1777
rect 27320 1743 27613 1777
rect 27647 1743 27949 1777
rect 27983 1743 28285 1777
rect 28319 1743 28621 1777
rect 28655 1743 28948 1777
rect 29000 1743 29293 1777
rect 29327 1743 29629 1777
rect 29663 1743 29965 1777
rect 29999 1743 30301 1777
rect 30335 1743 30628 1777
rect 30680 1743 30973 1777
rect 31007 1743 31309 1777
rect 31343 1743 31645 1777
rect 31679 1743 31981 1777
rect 32015 1743 32308 1777
rect 32360 1743 32653 1777
rect 32687 1743 32989 1777
rect 33023 1743 33325 1777
rect 33359 1743 33661 1777
rect 33695 1743 33988 1777
rect 34040 1743 34333 1777
rect 34367 1743 34669 1777
rect 34703 1743 35005 1777
rect 35039 1743 35341 1777
rect 35375 1743 35668 1777
rect 35720 1743 36013 1777
rect 36047 1743 36349 1777
rect 36383 1743 36685 1777
rect 36719 1743 37021 1777
rect 37055 1743 37348 1777
rect 37400 1743 37693 1777
rect 37727 1743 38029 1777
rect 38063 1743 38365 1777
rect 38399 1743 38701 1777
rect 38735 1743 39028 1777
rect 39080 1743 39373 1777
rect 39407 1743 39709 1777
rect 39743 1743 40045 1777
rect 40079 1743 40381 1777
rect 40415 1743 40708 1777
rect 40760 1743 41053 1777
rect 41087 1743 41852 1777
rect 2120 1734 3748 1743
rect 3800 1734 5428 1743
rect 5480 1734 7108 1743
rect 7160 1734 8788 1743
rect 8840 1734 10468 1743
rect 10520 1734 12148 1743
rect 12200 1734 13828 1743
rect 13880 1734 15508 1743
rect 15560 1734 17188 1743
rect 17240 1734 18868 1743
rect 18920 1734 20548 1743
rect 20600 1734 22228 1743
rect 22280 1734 23908 1743
rect 23960 1734 25588 1743
rect 25640 1734 27268 1743
rect 27320 1734 28948 1743
rect 29000 1734 30628 1743
rect 30680 1734 32308 1743
rect 32360 1734 33988 1743
rect 34040 1734 35668 1743
rect 35720 1734 37348 1743
rect 37400 1734 39028 1743
rect 39080 1734 40708 1743
rect 40760 1734 41852 1743
rect 1646 1648 41852 1734
<< via1 >>
rect 2068 31401 2120 31410
rect 3748 31401 3800 31410
rect 5428 31401 5480 31410
rect 7108 31401 7160 31410
rect 8788 31401 8840 31410
rect 10468 31401 10520 31410
rect 12148 31401 12200 31410
rect 13828 31401 13880 31410
rect 15508 31401 15560 31410
rect 17188 31401 17240 31410
rect 18868 31401 18920 31410
rect 20548 31401 20600 31410
rect 22228 31401 22280 31410
rect 23908 31401 23960 31410
rect 25588 31401 25640 31410
rect 27268 31401 27320 31410
rect 28948 31401 29000 31410
rect 30628 31401 30680 31410
rect 32308 31401 32360 31410
rect 33988 31401 34040 31410
rect 35668 31401 35720 31410
rect 37348 31401 37400 31410
rect 39028 31401 39080 31410
rect 40708 31401 40760 31410
rect 2068 31367 2077 31401
rect 2077 31367 2111 31401
rect 2111 31367 2120 31401
rect 3748 31367 3757 31401
rect 3757 31367 3791 31401
rect 3791 31367 3800 31401
rect 5428 31367 5437 31401
rect 5437 31367 5471 31401
rect 5471 31367 5480 31401
rect 7108 31367 7117 31401
rect 7117 31367 7151 31401
rect 7151 31367 7160 31401
rect 8788 31367 8797 31401
rect 8797 31367 8831 31401
rect 8831 31367 8840 31401
rect 10468 31367 10477 31401
rect 10477 31367 10511 31401
rect 10511 31367 10520 31401
rect 12148 31367 12157 31401
rect 12157 31367 12191 31401
rect 12191 31367 12200 31401
rect 13828 31367 13837 31401
rect 13837 31367 13871 31401
rect 13871 31367 13880 31401
rect 15508 31367 15517 31401
rect 15517 31367 15551 31401
rect 15551 31367 15560 31401
rect 17188 31367 17197 31401
rect 17197 31367 17231 31401
rect 17231 31367 17240 31401
rect 18868 31367 18877 31401
rect 18877 31367 18911 31401
rect 18911 31367 18920 31401
rect 20548 31367 20557 31401
rect 20557 31367 20591 31401
rect 20591 31367 20600 31401
rect 22228 31367 22237 31401
rect 22237 31367 22271 31401
rect 22271 31367 22280 31401
rect 23908 31367 23917 31401
rect 23917 31367 23951 31401
rect 23951 31367 23960 31401
rect 25588 31367 25597 31401
rect 25597 31367 25631 31401
rect 25631 31367 25640 31401
rect 27268 31367 27277 31401
rect 27277 31367 27311 31401
rect 27311 31367 27320 31401
rect 28948 31367 28957 31401
rect 28957 31367 28991 31401
rect 28991 31367 29000 31401
rect 30628 31367 30637 31401
rect 30637 31367 30671 31401
rect 30671 31367 30680 31401
rect 32308 31367 32317 31401
rect 32317 31367 32351 31401
rect 32351 31367 32360 31401
rect 33988 31367 33997 31401
rect 33997 31367 34031 31401
rect 34031 31367 34040 31401
rect 35668 31367 35677 31401
rect 35677 31367 35711 31401
rect 35711 31367 35720 31401
rect 37348 31367 37357 31401
rect 37357 31367 37391 31401
rect 37391 31367 37400 31401
rect 39028 31367 39037 31401
rect 39037 31367 39071 31401
rect 39071 31367 39080 31401
rect 40708 31367 40717 31401
rect 40717 31367 40751 31401
rect 40751 31367 40760 31401
rect 2068 31358 2120 31367
rect 3748 31358 3800 31367
rect 5428 31358 5480 31367
rect 7108 31358 7160 31367
rect 8788 31358 8840 31367
rect 10468 31358 10520 31367
rect 12148 31358 12200 31367
rect 13828 31358 13880 31367
rect 15508 31358 15560 31367
rect 17188 31358 17240 31367
rect 18868 31358 18920 31367
rect 20548 31358 20600 31367
rect 22228 31358 22280 31367
rect 23908 31358 23960 31367
rect 25588 31358 25640 31367
rect 27268 31358 27320 31367
rect 28948 31358 29000 31367
rect 30628 31358 30680 31367
rect 32308 31358 32360 31367
rect 33988 31358 34040 31367
rect 35668 31358 35720 31367
rect 37348 31358 37400 31367
rect 39028 31358 39080 31367
rect 40708 31358 40760 31367
rect 1732 31009 1784 31018
rect 1732 30975 1741 31009
rect 1741 30975 1775 31009
rect 1775 30975 1784 31009
rect 1732 30966 1784 30975
rect 41714 31009 41766 31018
rect 41714 30975 41723 31009
rect 41723 30975 41757 31009
rect 41757 30975 41766 31009
rect 41714 30966 41766 30975
rect 1732 30673 1784 30682
rect 1732 30639 1741 30673
rect 1741 30639 1775 30673
rect 1775 30639 1784 30673
rect 1732 30630 1784 30639
rect 41714 30673 41766 30682
rect 41714 30639 41723 30673
rect 41723 30639 41757 30673
rect 41757 30639 41766 30673
rect 41714 30630 41766 30639
rect 1732 30337 1784 30346
rect 1732 30303 1741 30337
rect 1741 30303 1775 30337
rect 1775 30303 1784 30337
rect 1732 30294 1784 30303
rect 41714 30337 41766 30346
rect 41714 30303 41723 30337
rect 41723 30303 41757 30337
rect 41757 30303 41766 30337
rect 41714 30294 41766 30303
rect 1732 30001 1784 30010
rect 1732 29967 1741 30001
rect 1741 29967 1775 30001
rect 1775 29967 1784 30001
rect 1732 29958 1784 29967
rect 41714 30001 41766 30010
rect 41714 29967 41723 30001
rect 41723 29967 41757 30001
rect 41757 29967 41766 30001
rect 41714 29958 41766 29967
rect 1732 29665 1784 29674
rect 1732 29631 1741 29665
rect 1741 29631 1775 29665
rect 1775 29631 1784 29665
rect 1732 29622 1784 29631
rect 41714 29665 41766 29674
rect 41714 29631 41723 29665
rect 41723 29631 41757 29665
rect 41757 29631 41766 29665
rect 41714 29622 41766 29631
rect 1732 29329 1784 29338
rect 1732 29295 1741 29329
rect 1741 29295 1775 29329
rect 1775 29295 1784 29329
rect 1732 29286 1784 29295
rect 41714 29329 41766 29338
rect 41714 29295 41723 29329
rect 41723 29295 41757 29329
rect 41757 29295 41766 29329
rect 41714 29286 41766 29295
rect 1732 28993 1784 29002
rect 1732 28959 1741 28993
rect 1741 28959 1775 28993
rect 1775 28959 1784 28993
rect 1732 28950 1784 28959
rect 41714 28993 41766 29002
rect 41714 28959 41723 28993
rect 41723 28959 41757 28993
rect 41757 28959 41766 28993
rect 41714 28950 41766 28959
rect 1732 28657 1784 28666
rect 1732 28623 1741 28657
rect 1741 28623 1775 28657
rect 1775 28623 1784 28657
rect 1732 28614 1784 28623
rect 41714 28657 41766 28666
rect 41714 28623 41723 28657
rect 41723 28623 41757 28657
rect 41757 28623 41766 28657
rect 41714 28614 41766 28623
rect 1732 28321 1784 28330
rect 1732 28287 1741 28321
rect 1741 28287 1775 28321
rect 1775 28287 1784 28321
rect 1732 28278 1784 28287
rect 41714 28321 41766 28330
rect 41714 28287 41723 28321
rect 41723 28287 41757 28321
rect 41757 28287 41766 28321
rect 41714 28278 41766 28287
rect 1732 27985 1784 27994
rect 1732 27951 1741 27985
rect 1741 27951 1775 27985
rect 1775 27951 1784 27985
rect 1732 27942 1784 27951
rect 41714 27985 41766 27994
rect 41714 27951 41723 27985
rect 41723 27951 41757 27985
rect 41757 27951 41766 27985
rect 41714 27942 41766 27951
rect 1732 27649 1784 27658
rect 1732 27615 1741 27649
rect 1741 27615 1775 27649
rect 1775 27615 1784 27649
rect 1732 27606 1784 27615
rect 41714 27649 41766 27658
rect 41714 27615 41723 27649
rect 41723 27615 41757 27649
rect 41757 27615 41766 27649
rect 41714 27606 41766 27615
rect 1732 27313 1784 27322
rect 1732 27279 1741 27313
rect 1741 27279 1775 27313
rect 1775 27279 1784 27313
rect 1732 27270 1784 27279
rect 41714 27313 41766 27322
rect 41714 27279 41723 27313
rect 41723 27279 41757 27313
rect 41757 27279 41766 27313
rect 41714 27270 41766 27279
rect 1732 26977 1784 26986
rect 1732 26943 1741 26977
rect 1741 26943 1775 26977
rect 1775 26943 1784 26977
rect 1732 26934 1784 26943
rect 41714 26977 41766 26986
rect 41714 26943 41723 26977
rect 41723 26943 41757 26977
rect 41757 26943 41766 26977
rect 41714 26934 41766 26943
rect 1732 26641 1784 26650
rect 1732 26607 1741 26641
rect 1741 26607 1775 26641
rect 1775 26607 1784 26641
rect 1732 26598 1784 26607
rect 41714 26641 41766 26650
rect 41714 26607 41723 26641
rect 41723 26607 41757 26641
rect 41757 26607 41766 26641
rect 41714 26598 41766 26607
rect 1732 26305 1784 26314
rect 1732 26271 1741 26305
rect 1741 26271 1775 26305
rect 1775 26271 1784 26305
rect 1732 26262 1784 26271
rect 41714 26305 41766 26314
rect 41714 26271 41723 26305
rect 41723 26271 41757 26305
rect 41757 26271 41766 26305
rect 41714 26262 41766 26271
rect 9941 26137 9993 26189
rect 1732 25969 1784 25978
rect 1732 25935 1741 25969
rect 1741 25935 1775 25969
rect 1775 25935 1784 25969
rect 1732 25926 1784 25935
rect 1732 25633 1784 25642
rect 1732 25599 1741 25633
rect 1741 25599 1775 25633
rect 1775 25599 1784 25633
rect 1732 25590 1784 25599
rect 1732 25297 1784 25306
rect 1732 25263 1741 25297
rect 1741 25263 1775 25297
rect 1775 25263 1784 25297
rect 1732 25254 1784 25263
rect 1732 24961 1784 24970
rect 1732 24927 1741 24961
rect 1741 24927 1775 24961
rect 1775 24927 1784 24961
rect 1732 24918 1784 24927
rect 1732 24625 1784 24634
rect 1732 24591 1741 24625
rect 1741 24591 1775 24625
rect 1775 24591 1784 24625
rect 1732 24582 1784 24591
rect 9861 24579 9913 24631
rect 1732 24289 1784 24298
rect 1732 24255 1741 24289
rect 1741 24255 1775 24289
rect 1775 24255 1784 24289
rect 1732 24246 1784 24255
rect 1732 23953 1784 23962
rect 1732 23919 1741 23953
rect 1741 23919 1775 23953
rect 1775 23919 1784 23953
rect 1732 23910 1784 23919
rect 1732 23617 1784 23626
rect 1732 23583 1741 23617
rect 1741 23583 1775 23617
rect 1775 23583 1784 23617
rect 1732 23574 1784 23583
rect 9781 23309 9833 23361
rect 1732 23281 1784 23290
rect 1732 23247 1741 23281
rect 1741 23247 1775 23281
rect 1775 23247 1784 23281
rect 1732 23238 1784 23247
rect 1732 22945 1784 22954
rect 1732 22911 1741 22945
rect 1741 22911 1775 22945
rect 1775 22911 1784 22945
rect 1732 22902 1784 22911
rect 1732 22609 1784 22618
rect 1732 22575 1741 22609
rect 1741 22575 1775 22609
rect 1775 22575 1784 22609
rect 1732 22566 1784 22575
rect 1732 22273 1784 22282
rect 1732 22239 1741 22273
rect 1741 22239 1775 22273
rect 1775 22239 1784 22273
rect 1732 22230 1784 22239
rect 1732 21937 1784 21946
rect 1732 21903 1741 21937
rect 1741 21903 1775 21937
rect 1775 21903 1784 21937
rect 1732 21894 1784 21903
rect 9701 21751 9753 21803
rect 1732 21601 1784 21610
rect 1732 21567 1741 21601
rect 1741 21567 1775 21601
rect 1775 21567 1784 21601
rect 1732 21558 1784 21567
rect 1732 21265 1784 21274
rect 1732 21231 1741 21265
rect 1741 21231 1775 21265
rect 1775 21231 1784 21265
rect 1732 21222 1784 21231
rect 1732 20929 1784 20938
rect 1732 20895 1741 20929
rect 1741 20895 1775 20929
rect 1775 20895 1784 20929
rect 1732 20886 1784 20895
rect 1732 20593 1784 20602
rect 1732 20559 1741 20593
rect 1741 20559 1775 20593
rect 1775 20559 1784 20593
rect 1732 20550 1784 20559
rect 1732 20257 1784 20266
rect 1732 20223 1741 20257
rect 1741 20223 1775 20257
rect 1775 20223 1784 20257
rect 1732 20214 1784 20223
rect 1732 19921 1784 19930
rect 1732 19887 1741 19921
rect 1741 19887 1775 19921
rect 1775 19887 1784 19921
rect 1732 19878 1784 19887
rect 1732 19585 1784 19594
rect 1732 19551 1741 19585
rect 1741 19551 1775 19585
rect 1775 19551 1784 19585
rect 1732 19542 1784 19551
rect 1732 19249 1784 19258
rect 1732 19215 1741 19249
rect 1741 19215 1775 19249
rect 1775 19215 1784 19249
rect 1732 19206 1784 19215
rect 1732 18913 1784 18922
rect 1732 18879 1741 18913
rect 1741 18879 1775 18913
rect 1775 18879 1784 18913
rect 1732 18870 1784 18879
rect 1732 18577 1784 18586
rect 1732 18543 1741 18577
rect 1741 18543 1775 18577
rect 1775 18543 1784 18577
rect 1732 18534 1784 18543
rect 1732 18241 1784 18250
rect 1732 18207 1741 18241
rect 1741 18207 1775 18241
rect 1775 18207 1784 18241
rect 1732 18198 1784 18207
rect 1732 17905 1784 17914
rect 1732 17871 1741 17905
rect 1741 17871 1775 17905
rect 1775 17871 1784 17905
rect 1732 17862 1784 17871
rect 1732 17569 1784 17578
rect 1732 17535 1741 17569
rect 1741 17535 1775 17569
rect 1775 17535 1784 17569
rect 1732 17526 1784 17535
rect 1732 17233 1784 17242
rect 1732 17199 1741 17233
rect 1741 17199 1775 17233
rect 1775 17199 1784 17233
rect 1732 17190 1784 17199
rect 1732 16897 1784 16906
rect 1732 16863 1741 16897
rect 1741 16863 1775 16897
rect 1775 16863 1784 16897
rect 1732 16854 1784 16863
rect 41714 25969 41766 25978
rect 41714 25935 41723 25969
rect 41723 25935 41757 25969
rect 41757 25935 41766 25969
rect 41714 25926 41766 25935
rect 41714 25633 41766 25642
rect 41714 25599 41723 25633
rect 41723 25599 41757 25633
rect 41757 25599 41766 25633
rect 41714 25590 41766 25599
rect 19408 25297 19460 25349
rect 20402 25297 20454 25349
rect 20656 25297 20708 25349
rect 21650 25297 21702 25349
rect 21904 25297 21956 25349
rect 22898 25297 22950 25349
rect 23152 25297 23204 25349
rect 24146 25297 24198 25349
rect 41714 25297 41766 25306
rect 41714 25263 41723 25297
rect 41723 25263 41757 25297
rect 41757 25263 41766 25297
rect 41714 25254 41766 25263
rect 41714 24961 41766 24970
rect 41714 24927 41723 24961
rect 41723 24927 41757 24961
rect 41757 24927 41766 24961
rect 41714 24918 41766 24927
rect 41714 24625 41766 24634
rect 41714 24591 41723 24625
rect 41723 24591 41757 24625
rect 41757 24591 41766 24625
rect 41714 24582 41766 24591
rect 41714 24289 41766 24298
rect 41714 24255 41723 24289
rect 41723 24255 41757 24289
rect 41757 24255 41766 24289
rect 41714 24246 41766 24255
rect 41714 23953 41766 23962
rect 41714 23919 41723 23953
rect 41723 23919 41757 23953
rect 41757 23919 41766 23953
rect 41714 23910 41766 23919
rect 41714 23617 41766 23626
rect 41714 23583 41723 23617
rect 41723 23583 41757 23617
rect 41757 23583 41766 23617
rect 41714 23574 41766 23583
rect 41714 23281 41766 23290
rect 41714 23247 41723 23281
rect 41723 23247 41757 23281
rect 41757 23247 41766 23281
rect 41714 23238 41766 23247
rect 41714 22945 41766 22954
rect 41714 22911 41723 22945
rect 41723 22911 41757 22945
rect 41757 22911 41766 22945
rect 41714 22902 41766 22911
rect 41714 22609 41766 22618
rect 41714 22575 41723 22609
rect 41723 22575 41757 22609
rect 41757 22575 41766 22609
rect 41714 22566 41766 22575
rect 41714 22273 41766 22282
rect 41714 22239 41723 22273
rect 41723 22239 41757 22273
rect 41757 22239 41766 22273
rect 41714 22230 41766 22239
rect 41714 21937 41766 21946
rect 41714 21903 41723 21937
rect 41723 21903 41757 21937
rect 41757 21903 41766 21937
rect 41714 21894 41766 21903
rect 41714 21601 41766 21610
rect 41714 21567 41723 21601
rect 41723 21567 41757 21601
rect 41757 21567 41766 21601
rect 41714 21558 41766 21567
rect 41714 21265 41766 21274
rect 41714 21231 41723 21265
rect 41723 21231 41757 21265
rect 41757 21231 41766 21265
rect 41714 21222 41766 21231
rect 41714 20929 41766 20938
rect 41714 20895 41723 20929
rect 41723 20895 41757 20929
rect 41757 20895 41766 20929
rect 41714 20886 41766 20895
rect 41714 20593 41766 20602
rect 41714 20559 41723 20593
rect 41723 20559 41757 20593
rect 41757 20559 41766 20593
rect 41714 20550 41766 20559
rect 41714 20257 41766 20266
rect 41714 20223 41723 20257
rect 41723 20223 41757 20257
rect 41757 20223 41766 20257
rect 41714 20214 41766 20223
rect 41714 19921 41766 19930
rect 41714 19887 41723 19921
rect 41723 19887 41757 19921
rect 41757 19887 41766 19921
rect 41714 19878 41766 19887
rect 41714 19585 41766 19594
rect 41714 19551 41723 19585
rect 41723 19551 41757 19585
rect 41757 19551 41766 19585
rect 41714 19542 41766 19551
rect 41714 19249 41766 19258
rect 41714 19215 41723 19249
rect 41723 19215 41757 19249
rect 41757 19215 41766 19249
rect 41714 19206 41766 19215
rect 41714 18913 41766 18922
rect 41714 18879 41723 18913
rect 41723 18879 41757 18913
rect 41757 18879 41766 18913
rect 41714 18870 41766 18879
rect 41714 18577 41766 18586
rect 41714 18543 41723 18577
rect 41723 18543 41757 18577
rect 41757 18543 41766 18577
rect 41714 18534 41766 18543
rect 41714 18241 41766 18250
rect 41714 18207 41723 18241
rect 41723 18207 41757 18241
rect 41757 18207 41766 18241
rect 41714 18198 41766 18207
rect 41714 17905 41766 17914
rect 41714 17871 41723 17905
rect 41723 17871 41757 17905
rect 41757 17871 41766 17905
rect 41714 17862 41766 17871
rect 41714 17569 41766 17578
rect 41714 17535 41723 17569
rect 41723 17535 41757 17569
rect 41757 17535 41766 17569
rect 41714 17526 41766 17535
rect 41714 17233 41766 17242
rect 41714 17199 41723 17233
rect 41723 17199 41757 17233
rect 41757 17199 41766 17233
rect 41714 17190 41766 17199
rect 41714 16897 41766 16906
rect 41714 16863 41723 16897
rect 41723 16863 41757 16897
rect 41757 16863 41766 16897
rect 41714 16854 41766 16863
rect 1732 16561 1784 16570
rect 1732 16527 1741 16561
rect 1741 16527 1775 16561
rect 1775 16527 1784 16561
rect 1732 16518 1784 16527
rect 1732 16225 1784 16234
rect 1732 16191 1741 16225
rect 1741 16191 1775 16225
rect 1775 16191 1784 16225
rect 1732 16182 1784 16191
rect 1732 15889 1784 15898
rect 1732 15855 1741 15889
rect 1741 15855 1775 15889
rect 1775 15855 1784 15889
rect 1732 15846 1784 15855
rect 1732 15553 1784 15562
rect 1732 15519 1741 15553
rect 1741 15519 1775 15553
rect 1775 15519 1784 15553
rect 1732 15510 1784 15519
rect 1732 15217 1784 15226
rect 1732 15183 1741 15217
rect 1741 15183 1775 15217
rect 1775 15183 1784 15217
rect 1732 15174 1784 15183
rect 1732 14881 1784 14890
rect 1732 14847 1741 14881
rect 1741 14847 1775 14881
rect 1775 14847 1784 14881
rect 1732 14838 1784 14847
rect 1732 14545 1784 14554
rect 1732 14511 1741 14545
rect 1741 14511 1775 14545
rect 1775 14511 1784 14545
rect 1732 14502 1784 14511
rect 1732 14209 1784 14218
rect 1732 14175 1741 14209
rect 1741 14175 1775 14209
rect 1775 14175 1784 14209
rect 1732 14166 1784 14175
rect 1732 13873 1784 13882
rect 1732 13839 1741 13873
rect 1741 13839 1775 13873
rect 1775 13839 1784 13873
rect 1732 13830 1784 13839
rect 1732 13537 1784 13546
rect 1732 13503 1741 13537
rect 1741 13503 1775 13537
rect 1775 13503 1784 13537
rect 1732 13494 1784 13503
rect 1732 13201 1784 13210
rect 1732 13167 1741 13201
rect 1741 13167 1775 13201
rect 1775 13167 1784 13201
rect 1732 13158 1784 13167
rect 1732 12865 1784 12874
rect 1732 12831 1741 12865
rect 1741 12831 1775 12865
rect 1775 12831 1784 12865
rect 1732 12822 1784 12831
rect 1732 12529 1784 12538
rect 1732 12495 1741 12529
rect 1741 12495 1775 12529
rect 1775 12495 1784 12529
rect 1732 12486 1784 12495
rect 1732 12193 1784 12202
rect 1732 12159 1741 12193
rect 1741 12159 1775 12193
rect 1775 12159 1784 12193
rect 1732 12150 1784 12159
rect 1732 11857 1784 11866
rect 1732 11823 1741 11857
rect 1741 11823 1775 11857
rect 1775 11823 1784 11857
rect 1732 11814 1784 11823
rect 1732 11521 1784 11530
rect 1732 11487 1741 11521
rect 1741 11487 1775 11521
rect 1775 11487 1784 11521
rect 1732 11478 1784 11487
rect 1732 11185 1784 11194
rect 1732 11151 1741 11185
rect 1741 11151 1775 11185
rect 1775 11151 1784 11185
rect 1732 11142 1784 11151
rect 1732 10849 1784 10858
rect 1732 10815 1741 10849
rect 1741 10815 1775 10849
rect 1775 10815 1784 10849
rect 1732 10806 1784 10815
rect 19408 10623 19460 10675
rect 20402 10623 20454 10675
rect 20656 10623 20708 10675
rect 21650 10623 21702 10675
rect 21904 10623 21956 10675
rect 22898 10623 22950 10675
rect 23152 10623 23204 10675
rect 24146 10623 24198 10675
rect 1732 10513 1784 10522
rect 1732 10479 1741 10513
rect 1741 10479 1775 10513
rect 1775 10479 1784 10513
rect 1732 10470 1784 10479
rect 1732 10177 1784 10186
rect 1732 10143 1741 10177
rect 1741 10143 1775 10177
rect 1775 10143 1784 10177
rect 1732 10134 1784 10143
rect 1732 9841 1784 9850
rect 1732 9807 1741 9841
rect 1741 9807 1775 9841
rect 1775 9807 1784 9841
rect 1732 9798 1784 9807
rect 41714 16561 41766 16570
rect 41714 16527 41723 16561
rect 41723 16527 41757 16561
rect 41757 16527 41766 16561
rect 41714 16518 41766 16527
rect 41714 16225 41766 16234
rect 41714 16191 41723 16225
rect 41723 16191 41757 16225
rect 41757 16191 41766 16225
rect 41714 16182 41766 16191
rect 41714 15889 41766 15898
rect 41714 15855 41723 15889
rect 41723 15855 41757 15889
rect 41757 15855 41766 15889
rect 41714 15846 41766 15855
rect 41714 15553 41766 15562
rect 41714 15519 41723 15553
rect 41723 15519 41757 15553
rect 41757 15519 41766 15553
rect 41714 15510 41766 15519
rect 41714 15217 41766 15226
rect 41714 15183 41723 15217
rect 41723 15183 41757 15217
rect 41757 15183 41766 15217
rect 41714 15174 41766 15183
rect 41714 14881 41766 14890
rect 41714 14847 41723 14881
rect 41723 14847 41757 14881
rect 41757 14847 41766 14881
rect 41714 14838 41766 14847
rect 41714 14545 41766 14554
rect 41714 14511 41723 14545
rect 41723 14511 41757 14545
rect 41757 14511 41766 14545
rect 41714 14502 41766 14511
rect 33853 14165 33905 14217
rect 41714 14209 41766 14218
rect 41714 14175 41723 14209
rect 41723 14175 41757 14209
rect 41757 14175 41766 14209
rect 41714 14166 41766 14175
rect 41714 13873 41766 13882
rect 41714 13839 41723 13873
rect 41723 13839 41757 13873
rect 41757 13839 41766 13873
rect 41714 13830 41766 13839
rect 41714 13537 41766 13546
rect 41714 13503 41723 13537
rect 41723 13503 41757 13537
rect 41757 13503 41766 13537
rect 41714 13494 41766 13503
rect 41714 13201 41766 13210
rect 41714 13167 41723 13201
rect 41723 13167 41757 13201
rect 41757 13167 41766 13201
rect 41714 13158 41766 13167
rect 41714 12865 41766 12874
rect 41714 12831 41723 12865
rect 41723 12831 41757 12865
rect 41757 12831 41766 12865
rect 41714 12822 41766 12831
rect 33773 12607 33825 12659
rect 41714 12529 41766 12538
rect 41714 12495 41723 12529
rect 41723 12495 41757 12529
rect 41757 12495 41766 12529
rect 41714 12486 41766 12495
rect 41714 12193 41766 12202
rect 41714 12159 41723 12193
rect 41723 12159 41757 12193
rect 41757 12159 41766 12193
rect 41714 12150 41766 12159
rect 41714 11857 41766 11866
rect 41714 11823 41723 11857
rect 41723 11823 41757 11857
rect 41757 11823 41766 11857
rect 41714 11814 41766 11823
rect 41714 11521 41766 11530
rect 41714 11487 41723 11521
rect 41723 11487 41757 11521
rect 41757 11487 41766 11521
rect 41714 11478 41766 11487
rect 33693 11337 33745 11389
rect 41714 11185 41766 11194
rect 41714 11151 41723 11185
rect 41723 11151 41757 11185
rect 41757 11151 41766 11185
rect 41714 11142 41766 11151
rect 41714 10849 41766 10858
rect 41714 10815 41723 10849
rect 41723 10815 41757 10849
rect 41757 10815 41766 10849
rect 41714 10806 41766 10815
rect 41714 10513 41766 10522
rect 41714 10479 41723 10513
rect 41723 10479 41757 10513
rect 41757 10479 41766 10513
rect 41714 10470 41766 10479
rect 41714 10177 41766 10186
rect 41714 10143 41723 10177
rect 41723 10143 41757 10177
rect 41757 10143 41766 10177
rect 41714 10134 41766 10143
rect 33613 9779 33665 9831
rect 41714 9841 41766 9850
rect 41714 9807 41723 9841
rect 41723 9807 41757 9841
rect 41757 9807 41766 9841
rect 41714 9798 41766 9807
rect 1732 9505 1784 9514
rect 1732 9471 1741 9505
rect 1741 9471 1775 9505
rect 1775 9471 1784 9505
rect 1732 9462 1784 9471
rect 41714 9505 41766 9514
rect 41714 9471 41723 9505
rect 41723 9471 41757 9505
rect 41757 9471 41766 9505
rect 41714 9462 41766 9471
rect 1732 9169 1784 9178
rect 1732 9135 1741 9169
rect 1741 9135 1775 9169
rect 1775 9135 1784 9169
rect 1732 9126 1784 9135
rect 41714 9169 41766 9178
rect 41714 9135 41723 9169
rect 41723 9135 41757 9169
rect 41757 9135 41766 9169
rect 41714 9126 41766 9135
rect 1732 8833 1784 8842
rect 1732 8799 1741 8833
rect 1741 8799 1775 8833
rect 1775 8799 1784 8833
rect 1732 8790 1784 8799
rect 41714 8833 41766 8842
rect 41714 8799 41723 8833
rect 41723 8799 41757 8833
rect 41757 8799 41766 8833
rect 41714 8790 41766 8799
rect 1732 8497 1784 8506
rect 1732 8463 1741 8497
rect 1741 8463 1775 8497
rect 1775 8463 1784 8497
rect 1732 8454 1784 8463
rect 41714 8497 41766 8506
rect 41714 8463 41723 8497
rect 41723 8463 41757 8497
rect 41757 8463 41766 8497
rect 41714 8454 41766 8463
rect 1732 8161 1784 8170
rect 1732 8127 1741 8161
rect 1741 8127 1775 8161
rect 1775 8127 1784 8161
rect 1732 8118 1784 8127
rect 41714 8161 41766 8170
rect 41714 8127 41723 8161
rect 41723 8127 41757 8161
rect 41757 8127 41766 8161
rect 41714 8118 41766 8127
rect 1732 7825 1784 7834
rect 1732 7791 1741 7825
rect 1741 7791 1775 7825
rect 1775 7791 1784 7825
rect 1732 7782 1784 7791
rect 41714 7825 41766 7834
rect 41714 7791 41723 7825
rect 41723 7791 41757 7825
rect 41757 7791 41766 7825
rect 41714 7782 41766 7791
rect 1732 7489 1784 7498
rect 1732 7455 1741 7489
rect 1741 7455 1775 7489
rect 1775 7455 1784 7489
rect 1732 7446 1784 7455
rect 41714 7489 41766 7498
rect 41714 7455 41723 7489
rect 41723 7455 41757 7489
rect 41757 7455 41766 7489
rect 41714 7446 41766 7455
rect 1732 7153 1784 7162
rect 1732 7119 1741 7153
rect 1741 7119 1775 7153
rect 1775 7119 1784 7153
rect 1732 7110 1784 7119
rect 41714 7153 41766 7162
rect 41714 7119 41723 7153
rect 41723 7119 41757 7153
rect 41757 7119 41766 7153
rect 41714 7110 41766 7119
rect 1732 6817 1784 6826
rect 1732 6783 1741 6817
rect 1741 6783 1775 6817
rect 1775 6783 1784 6817
rect 1732 6774 1784 6783
rect 41714 6817 41766 6826
rect 41714 6783 41723 6817
rect 41723 6783 41757 6817
rect 41757 6783 41766 6817
rect 41714 6774 41766 6783
rect 1732 6481 1784 6490
rect 1732 6447 1741 6481
rect 1741 6447 1775 6481
rect 1775 6447 1784 6481
rect 1732 6438 1784 6447
rect 41714 6481 41766 6490
rect 41714 6447 41723 6481
rect 41723 6447 41757 6481
rect 41757 6447 41766 6481
rect 41714 6438 41766 6447
rect 1732 6145 1784 6154
rect 1732 6111 1741 6145
rect 1741 6111 1775 6145
rect 1775 6111 1784 6145
rect 1732 6102 1784 6111
rect 41714 6145 41766 6154
rect 41714 6111 41723 6145
rect 41723 6111 41757 6145
rect 41757 6111 41766 6145
rect 41714 6102 41766 6111
rect 1732 5809 1784 5818
rect 1732 5775 1741 5809
rect 1741 5775 1775 5809
rect 1775 5775 1784 5809
rect 1732 5766 1784 5775
rect 41714 5809 41766 5818
rect 41714 5775 41723 5809
rect 41723 5775 41757 5809
rect 41757 5775 41766 5809
rect 41714 5766 41766 5775
rect 1732 5473 1784 5482
rect 1732 5439 1741 5473
rect 1741 5439 1775 5473
rect 1775 5439 1784 5473
rect 1732 5430 1784 5439
rect 41714 5473 41766 5482
rect 41714 5439 41723 5473
rect 41723 5439 41757 5473
rect 41757 5439 41766 5473
rect 41714 5430 41766 5439
rect 1732 5137 1784 5146
rect 1732 5103 1741 5137
rect 1741 5103 1775 5137
rect 1775 5103 1784 5137
rect 1732 5094 1784 5103
rect 41714 5137 41766 5146
rect 41714 5103 41723 5137
rect 41723 5103 41757 5137
rect 41757 5103 41766 5137
rect 41714 5094 41766 5103
rect 1732 4801 1784 4810
rect 1732 4767 1741 4801
rect 1741 4767 1775 4801
rect 1775 4767 1784 4801
rect 1732 4758 1784 4767
rect 41714 4801 41766 4810
rect 41714 4767 41723 4801
rect 41723 4767 41757 4801
rect 41757 4767 41766 4801
rect 41714 4758 41766 4767
rect 1732 4465 1784 4474
rect 1732 4431 1741 4465
rect 1741 4431 1775 4465
rect 1775 4431 1784 4465
rect 1732 4422 1784 4431
rect 41714 4465 41766 4474
rect 41714 4431 41723 4465
rect 41723 4431 41757 4465
rect 41757 4431 41766 4465
rect 41714 4422 41766 4431
rect 1732 4129 1784 4138
rect 1732 4095 1741 4129
rect 1741 4095 1775 4129
rect 1775 4095 1784 4129
rect 1732 4086 1784 4095
rect 41714 4129 41766 4138
rect 41714 4095 41723 4129
rect 41723 4095 41757 4129
rect 41757 4095 41766 4129
rect 41714 4086 41766 4095
rect 1732 3793 1784 3802
rect 1732 3759 1741 3793
rect 1741 3759 1775 3793
rect 1775 3759 1784 3793
rect 1732 3750 1784 3759
rect 41714 3793 41766 3802
rect 41714 3759 41723 3793
rect 41723 3759 41757 3793
rect 41757 3759 41766 3793
rect 41714 3750 41766 3759
rect 1732 3457 1784 3466
rect 1732 3423 1741 3457
rect 1741 3423 1775 3457
rect 1775 3423 1784 3457
rect 1732 3414 1784 3423
rect 41714 3457 41766 3466
rect 41714 3423 41723 3457
rect 41723 3423 41757 3457
rect 41757 3423 41766 3457
rect 41714 3414 41766 3423
rect 1732 3121 1784 3130
rect 1732 3087 1741 3121
rect 1741 3087 1775 3121
rect 1775 3087 1784 3121
rect 1732 3078 1784 3087
rect 41714 3121 41766 3130
rect 41714 3087 41723 3121
rect 41723 3087 41757 3121
rect 41757 3087 41766 3121
rect 41714 3078 41766 3087
rect 1732 2785 1784 2794
rect 1732 2751 1741 2785
rect 1741 2751 1775 2785
rect 1775 2751 1784 2785
rect 1732 2742 1784 2751
rect 41714 2785 41766 2794
rect 41714 2751 41723 2785
rect 41723 2751 41757 2785
rect 41757 2751 41766 2785
rect 41714 2742 41766 2751
rect 1732 2449 1784 2458
rect 1732 2415 1741 2449
rect 1741 2415 1775 2449
rect 1775 2415 1784 2449
rect 1732 2406 1784 2415
rect 41714 2449 41766 2458
rect 41714 2415 41723 2449
rect 41723 2415 41757 2449
rect 41757 2415 41766 2449
rect 41714 2406 41766 2415
rect 1732 2113 1784 2122
rect 1732 2079 1741 2113
rect 1741 2079 1775 2113
rect 1775 2079 1784 2113
rect 1732 2070 1784 2079
rect 41714 2113 41766 2122
rect 41714 2079 41723 2113
rect 41723 2079 41757 2113
rect 41757 2079 41766 2113
rect 41714 2070 41766 2079
rect 2068 1777 2120 1786
rect 3748 1777 3800 1786
rect 5428 1777 5480 1786
rect 7108 1777 7160 1786
rect 8788 1777 8840 1786
rect 10468 1777 10520 1786
rect 12148 1777 12200 1786
rect 13828 1777 13880 1786
rect 15508 1777 15560 1786
rect 17188 1777 17240 1786
rect 18868 1777 18920 1786
rect 20548 1777 20600 1786
rect 22228 1777 22280 1786
rect 23908 1777 23960 1786
rect 25588 1777 25640 1786
rect 27268 1777 27320 1786
rect 28948 1777 29000 1786
rect 30628 1777 30680 1786
rect 32308 1777 32360 1786
rect 33988 1777 34040 1786
rect 35668 1777 35720 1786
rect 37348 1777 37400 1786
rect 39028 1777 39080 1786
rect 40708 1777 40760 1786
rect 2068 1743 2077 1777
rect 2077 1743 2111 1777
rect 2111 1743 2120 1777
rect 3748 1743 3757 1777
rect 3757 1743 3791 1777
rect 3791 1743 3800 1777
rect 5428 1743 5437 1777
rect 5437 1743 5471 1777
rect 5471 1743 5480 1777
rect 7108 1743 7117 1777
rect 7117 1743 7151 1777
rect 7151 1743 7160 1777
rect 8788 1743 8797 1777
rect 8797 1743 8831 1777
rect 8831 1743 8840 1777
rect 10468 1743 10477 1777
rect 10477 1743 10511 1777
rect 10511 1743 10520 1777
rect 12148 1743 12157 1777
rect 12157 1743 12191 1777
rect 12191 1743 12200 1777
rect 13828 1743 13837 1777
rect 13837 1743 13871 1777
rect 13871 1743 13880 1777
rect 15508 1743 15517 1777
rect 15517 1743 15551 1777
rect 15551 1743 15560 1777
rect 17188 1743 17197 1777
rect 17197 1743 17231 1777
rect 17231 1743 17240 1777
rect 18868 1743 18877 1777
rect 18877 1743 18911 1777
rect 18911 1743 18920 1777
rect 20548 1743 20557 1777
rect 20557 1743 20591 1777
rect 20591 1743 20600 1777
rect 22228 1743 22237 1777
rect 22237 1743 22271 1777
rect 22271 1743 22280 1777
rect 23908 1743 23917 1777
rect 23917 1743 23951 1777
rect 23951 1743 23960 1777
rect 25588 1743 25597 1777
rect 25597 1743 25631 1777
rect 25631 1743 25640 1777
rect 27268 1743 27277 1777
rect 27277 1743 27311 1777
rect 27311 1743 27320 1777
rect 28948 1743 28957 1777
rect 28957 1743 28991 1777
rect 28991 1743 29000 1777
rect 30628 1743 30637 1777
rect 30637 1743 30671 1777
rect 30671 1743 30680 1777
rect 32308 1743 32317 1777
rect 32317 1743 32351 1777
rect 32351 1743 32360 1777
rect 33988 1743 33997 1777
rect 33997 1743 34031 1777
rect 34031 1743 34040 1777
rect 35668 1743 35677 1777
rect 35677 1743 35711 1777
rect 35711 1743 35720 1777
rect 37348 1743 37357 1777
rect 37357 1743 37391 1777
rect 37391 1743 37400 1777
rect 39028 1743 39037 1777
rect 39037 1743 39071 1777
rect 39071 1743 39080 1777
rect 40708 1743 40717 1777
rect 40717 1743 40751 1777
rect 40751 1743 40760 1777
rect 2068 1734 2120 1743
rect 3748 1734 3800 1743
rect 5428 1734 5480 1743
rect 7108 1734 7160 1743
rect 8788 1734 8840 1743
rect 10468 1734 10520 1743
rect 12148 1734 12200 1743
rect 13828 1734 13880 1743
rect 15508 1734 15560 1743
rect 17188 1734 17240 1743
rect 18868 1734 18920 1743
rect 20548 1734 20600 1743
rect 22228 1734 22280 1743
rect 23908 1734 23960 1743
rect 25588 1734 25640 1743
rect 27268 1734 27320 1743
rect 28948 1734 29000 1743
rect 30628 1734 30680 1743
rect 32308 1734 32360 1743
rect 33988 1734 34040 1743
rect 35668 1734 35720 1743
rect 37348 1734 37400 1743
rect 39028 1734 39080 1743
rect 40708 1734 40760 1743
<< metal2 >>
rect 1646 31018 1870 31496
rect 2066 31412 2122 31421
rect 2066 31347 2122 31356
rect 3746 31412 3802 31421
rect 3746 31347 3802 31356
rect 5426 31412 5482 31421
rect 5426 31347 5482 31356
rect 7106 31412 7162 31421
rect 7106 31347 7162 31356
rect 8786 31412 8842 31421
rect 8786 31347 8842 31356
rect 10466 31412 10522 31421
rect 10466 31347 10522 31356
rect 12146 31412 12202 31421
rect 12146 31347 12202 31356
rect 13826 31412 13882 31421
rect 13826 31347 13882 31356
rect 15506 31412 15562 31421
rect 15506 31347 15562 31356
rect 17186 31412 17242 31421
rect 17186 31347 17242 31356
rect 18866 31412 18922 31421
rect 18866 31347 18922 31356
rect 20546 31412 20602 31421
rect 20546 31347 20602 31356
rect 22226 31412 22282 31421
rect 22226 31347 22282 31356
rect 23906 31412 23962 31421
rect 23906 31347 23962 31356
rect 25586 31412 25642 31421
rect 25586 31347 25642 31356
rect 27266 31412 27322 31421
rect 27266 31347 27322 31356
rect 28946 31412 29002 31421
rect 28946 31347 29002 31356
rect 30626 31412 30682 31421
rect 30626 31347 30682 31356
rect 32306 31412 32362 31421
rect 32306 31347 32362 31356
rect 33986 31412 34042 31421
rect 33986 31347 34042 31356
rect 35666 31412 35722 31421
rect 35666 31347 35722 31356
rect 37346 31412 37402 31421
rect 37346 31347 37402 31356
rect 39026 31412 39082 31421
rect 39026 31347 39082 31356
rect 40706 31412 40762 31421
rect 40706 31347 40762 31356
rect 1646 30966 1732 31018
rect 1784 30966 1870 31018
rect 1646 30684 1870 30966
rect 1646 30628 1730 30684
rect 1786 30628 1870 30684
rect 1646 30346 1870 30628
rect 1646 30294 1732 30346
rect 1784 30294 1870 30346
rect 1646 30010 1870 30294
rect 41628 31018 41852 31496
rect 41628 30966 41714 31018
rect 41766 30966 41852 31018
rect 41628 30684 41852 30966
rect 41628 30628 41712 30684
rect 41768 30628 41852 30684
rect 41628 30346 41852 30628
rect 41628 30294 41714 30346
rect 41766 30294 41852 30346
rect 1646 29958 1732 30010
rect 1784 29958 1870 30010
rect 1646 29674 1870 29958
rect 40584 30008 40640 30017
rect 40584 29943 40640 29952
rect 41628 30010 41852 30294
rect 41628 29958 41714 30010
rect 41766 29958 41852 30010
rect 37447 29903 37503 29912
rect 1646 29622 1732 29674
rect 1784 29622 1870 29674
rect 1646 29338 1870 29622
rect 1646 29286 1732 29338
rect 1784 29286 1870 29338
rect 1646 29004 1870 29286
rect 1646 28948 1730 29004
rect 1786 28948 1870 29004
rect 1646 28666 1870 28948
rect 1646 28614 1732 28666
rect 1784 28614 1870 28666
rect 1646 28330 1870 28614
rect 1646 28278 1732 28330
rect 1784 28278 1870 28330
rect 1646 27994 1870 28278
rect 1646 27942 1732 27994
rect 1784 27942 1870 27994
rect 1646 27658 1870 27942
rect 1646 27606 1732 27658
rect 1784 27606 1870 27658
rect 1646 27324 1870 27606
rect 1646 27268 1730 27324
rect 1786 27268 1870 27324
rect 1646 26986 1870 27268
rect 1646 26934 1732 26986
rect 1784 26934 1870 26986
rect 1646 26650 1870 26934
rect 1646 26598 1732 26650
rect 1784 26598 1870 26650
rect 1646 26314 1870 26598
rect 1646 26262 1732 26314
rect 1784 26262 1870 26314
rect 34066 29823 34164 29851
rect 37447 29838 37503 29847
rect 1646 25978 1870 26262
rect 8500 26262 8556 26271
rect 8500 26197 8556 26206
rect 9445 26191 9501 26200
rect 9445 26126 9501 26135
rect 9939 26191 9995 26200
rect 9939 26126 9995 26135
rect 1646 25926 1732 25978
rect 1784 25926 1870 25978
rect 1646 25644 1870 25926
rect 1646 25588 1730 25644
rect 1786 25588 1870 25644
rect 1646 25306 1870 25588
rect 25969 25607 26025 25616
rect 25969 25542 26025 25551
rect 25983 25520 26011 25542
rect 1646 25254 1732 25306
rect 1784 25254 1870 25306
rect 19406 25351 19462 25360
rect 19406 25286 19462 25295
rect 20400 25351 20456 25360
rect 20400 25286 20456 25295
rect 20654 25351 20710 25360
rect 20654 25286 20710 25295
rect 21648 25351 21704 25360
rect 21648 25286 21704 25295
rect 21902 25351 21958 25360
rect 21902 25286 21958 25295
rect 22896 25351 22952 25360
rect 22896 25286 22952 25295
rect 23150 25351 23206 25360
rect 23150 25286 23206 25295
rect 24144 25351 24200 25360
rect 24144 25286 24200 25295
rect 1646 24970 1870 25254
rect 1646 24918 1732 24970
rect 1784 24918 1870 24970
rect 1646 24634 1870 24918
rect 1646 24582 1732 24634
rect 1784 24582 1870 24634
rect 1646 24298 1870 24582
rect 9445 24633 9501 24642
rect 8500 24562 8556 24571
rect 9445 24568 9501 24577
rect 9859 24633 9915 24642
rect 9859 24568 9915 24577
rect 8500 24497 8556 24506
rect 1646 24246 1732 24298
rect 1784 24246 1870 24298
rect 26107 24255 26135 25548
rect 1646 23964 1870 24246
rect 26093 24246 26149 24255
rect 26093 24181 26149 24190
rect 1646 23908 1730 23964
rect 1786 23908 1870 23964
rect 1646 23626 1870 23908
rect 1646 23574 1732 23626
rect 1784 23574 1870 23626
rect 1646 23290 1870 23574
rect 8500 23434 8556 23443
rect 8500 23369 8556 23378
rect 9445 23363 9501 23372
rect 9445 23298 9501 23307
rect 9779 23363 9835 23372
rect 9779 23298 9835 23307
rect 1646 23238 1732 23290
rect 1784 23238 1870 23290
rect 1646 22954 1870 23238
rect 1646 22902 1732 22954
rect 1784 22902 1870 22954
rect 1646 22618 1870 22902
rect 27902 22795 27958 22804
rect 27902 22730 27958 22739
rect 1646 22566 1732 22618
rect 1784 22566 1870 22618
rect 1646 22284 1870 22566
rect 1646 22228 1730 22284
rect 1786 22228 1870 22284
rect 1646 21946 1870 22228
rect 1646 21894 1732 21946
rect 1784 21894 1870 21946
rect 1646 21610 1870 21894
rect 9445 21805 9501 21814
rect 8500 21734 8556 21743
rect 9445 21740 9501 21749
rect 9699 21805 9755 21814
rect 9699 21740 9755 21749
rect 8500 21669 8556 21678
rect 1646 21558 1732 21610
rect 1784 21558 1870 21610
rect 1646 21274 1870 21558
rect 9582 21478 9638 21487
rect 27916 21445 27944 22730
rect 9582 21413 9638 21422
rect 1646 21222 1732 21274
rect 1784 21222 1870 21274
rect 1646 20938 1870 21222
rect 1646 20886 1732 20938
rect 1784 20886 1870 20938
rect 1646 20604 1870 20886
rect 1646 20548 1730 20604
rect 1786 20548 1870 20604
rect 1646 20266 1870 20548
rect 2645 20341 2701 20350
rect 2645 20276 2701 20285
rect 1646 20214 1732 20266
rect 1784 20214 1870 20266
rect 1646 19930 1870 20214
rect 1646 19878 1732 19930
rect 1784 19878 1870 19930
rect 1646 19594 1870 19878
rect 1646 19542 1732 19594
rect 1784 19542 1870 19594
rect 1646 19258 1870 19542
rect 1646 19206 1732 19258
rect 1784 19206 1870 19258
rect 1646 18924 1870 19206
rect 1646 18868 1730 18924
rect 1786 18868 1870 18924
rect 1646 18586 1870 18868
rect 1646 18534 1732 18586
rect 1784 18534 1870 18586
rect 1646 18250 1870 18534
rect 1646 18198 1732 18250
rect 1784 18198 1870 18250
rect 1646 17914 1870 18198
rect 1646 17862 1732 17914
rect 1784 17862 1870 17914
rect 1646 17578 1870 17862
rect 1646 17526 1732 17578
rect 1784 17526 1870 17578
rect 1646 17244 1870 17526
rect 1646 17188 1730 17244
rect 1786 17188 1870 17244
rect 1646 16906 1870 17188
rect 1646 16854 1732 16906
rect 1784 16854 1870 16906
rect 1646 16570 1870 16854
rect 1646 16518 1732 16570
rect 1784 16518 1870 16570
rect 1646 16234 1870 16518
rect 1646 16182 1732 16234
rect 1784 16182 1870 16234
rect 1646 15898 1870 16182
rect 1646 15846 1732 15898
rect 1784 15846 1870 15898
rect 1646 15564 1870 15846
rect 1646 15508 1730 15564
rect 1786 15508 1870 15564
rect 1646 15226 1870 15508
rect 1646 15174 1732 15226
rect 1784 15174 1870 15226
rect 1646 14890 1870 15174
rect 1646 14838 1732 14890
rect 1784 14838 1870 14890
rect 1646 14554 1870 14838
rect 1646 14502 1732 14554
rect 1784 14502 1870 14554
rect 1646 14218 1870 14502
rect 1646 14166 1732 14218
rect 1784 14166 1870 14218
rect 1646 13884 1870 14166
rect 1646 13828 1730 13884
rect 1786 13828 1870 13884
rect 1646 13546 1870 13828
rect 1646 13494 1732 13546
rect 1784 13494 1870 13546
rect 1646 13210 1870 13494
rect 1646 13158 1732 13210
rect 1784 13158 1870 13210
rect 9498 13233 9554 13242
rect 9498 13168 9554 13177
rect 1646 12874 1870 13158
rect 1646 12822 1732 12874
rect 1784 12822 1870 12874
rect 1646 12538 1870 12822
rect 1646 12486 1732 12538
rect 1784 12486 1870 12538
rect 1646 12204 1870 12486
rect 1646 12148 1730 12204
rect 1786 12148 1870 12204
rect 1646 11866 1870 12148
rect 1646 11814 1732 11866
rect 1784 11814 1870 11866
rect 1646 11530 1870 11814
rect 1646 11478 1732 11530
rect 1784 11478 1870 11530
rect 1646 11194 1870 11478
rect 1646 11142 1732 11194
rect 1784 11142 1870 11194
rect 1646 10858 1870 11142
rect 1646 10806 1732 10858
rect 1784 10806 1870 10858
rect 1646 10524 1870 10806
rect 1646 10468 1730 10524
rect 1786 10468 1870 10524
rect 1646 10186 1870 10468
rect 9498 10442 9554 10451
rect 9498 10377 9554 10386
rect 1646 10134 1732 10186
rect 1784 10134 1870 10186
rect 1646 9850 1870 10134
rect 1646 9798 1732 9850
rect 1784 9798 1870 9850
rect 1646 9514 1870 9798
rect 1646 9462 1732 9514
rect 1784 9462 1870 9514
rect 1646 9178 1870 9462
rect 1646 9126 1732 9178
rect 1784 9126 1870 9178
rect 1646 8844 1870 9126
rect 9498 8991 9554 9000
rect 9498 8926 9554 8935
rect 1646 8788 1730 8844
rect 1786 8788 1870 8844
rect 1646 8506 1870 8788
rect 1646 8454 1732 8506
rect 1784 8454 1870 8506
rect 1646 8170 1870 8454
rect 1646 8118 1732 8170
rect 1784 8118 1870 8170
rect 1646 7834 1870 8118
rect 1646 7782 1732 7834
rect 1784 7782 1870 7834
rect 1646 7498 1870 7782
rect 9498 7593 9554 7602
rect 9498 7528 9554 7537
rect 1646 7446 1732 7498
rect 1784 7446 1870 7498
rect 1646 7164 1870 7446
rect 1646 7108 1730 7164
rect 1786 7108 1870 7164
rect 1646 6826 1870 7108
rect 1646 6774 1732 6826
rect 1784 6774 1870 6826
rect 1646 6490 1870 6774
rect 1646 6438 1732 6490
rect 1784 6438 1870 6490
rect 1646 6154 1870 6438
rect 1646 6102 1732 6154
rect 1784 6102 1870 6154
rect 1646 5818 1870 6102
rect 1646 5766 1732 5818
rect 1784 5766 1870 5818
rect 1646 5484 1870 5766
rect 1646 5428 1730 5484
rect 1786 5428 1870 5484
rect 1646 5146 1870 5428
rect 1646 5094 1732 5146
rect 1784 5094 1870 5146
rect 1646 4810 1870 5094
rect 2858 4892 2914 4901
rect 2858 4827 2914 4836
rect 1646 4758 1732 4810
rect 1784 4758 1870 4810
rect 1646 4474 1870 4758
rect 1646 4422 1732 4474
rect 1784 4422 1870 4474
rect 1646 4138 1870 4422
rect 1646 4086 1732 4138
rect 1784 4086 1870 4138
rect 1646 3804 1870 4086
rect 1646 3748 1730 3804
rect 1786 3748 1870 3804
rect 1646 3466 1870 3748
rect 1646 3414 1732 3466
rect 1784 3414 1870 3466
rect 1646 3130 1870 3414
rect 9596 3321 9624 21413
rect 34066 14555 34094 29823
rect 41628 29674 41852 29958
rect 41628 29622 41714 29674
rect 41766 29622 41852 29674
rect 41628 29338 41852 29622
rect 41628 29286 41714 29338
rect 41766 29286 41852 29338
rect 41628 29004 41852 29286
rect 41628 28948 41712 29004
rect 41768 28948 41852 29004
rect 41628 28666 41852 28948
rect 41628 28614 41714 28666
rect 41766 28614 41852 28666
rect 41628 28330 41852 28614
rect 41628 28278 41714 28330
rect 41766 28278 41852 28330
rect 41628 27994 41852 28278
rect 41628 27942 41714 27994
rect 41766 27942 41852 27994
rect 41628 27658 41852 27942
rect 41628 27606 41714 27658
rect 41766 27606 41852 27658
rect 41628 27324 41852 27606
rect 41628 27268 41712 27324
rect 41768 27268 41852 27324
rect 41628 26986 41852 27268
rect 41628 26934 41714 26986
rect 41766 26934 41852 26986
rect 41628 26650 41852 26934
rect 41628 26598 41714 26650
rect 41766 26598 41852 26650
rect 41628 26314 41852 26598
rect 41628 26262 41714 26314
rect 41766 26262 41852 26314
rect 41628 25978 41852 26262
rect 41628 25926 41714 25978
rect 41766 25926 41852 25978
rect 41628 25644 41852 25926
rect 34136 25607 34192 25616
rect 34136 25542 34192 25551
rect 41628 25588 41712 25644
rect 41768 25588 41852 25644
rect 41628 25306 41852 25588
rect 41628 25254 41714 25306
rect 41766 25254 41852 25306
rect 41628 24970 41852 25254
rect 41628 24918 41714 24970
rect 41766 24918 41852 24970
rect 41628 24634 41852 24918
rect 41628 24582 41714 24634
rect 41766 24582 41852 24634
rect 41628 24298 41852 24582
rect 34136 24246 34192 24255
rect 34136 24181 34192 24190
rect 41628 24246 41714 24298
rect 41766 24246 41852 24298
rect 41628 23964 41852 24246
rect 41628 23908 41712 23964
rect 41768 23908 41852 23964
rect 41628 23626 41852 23908
rect 41628 23574 41714 23626
rect 41766 23574 41852 23626
rect 41628 23290 41852 23574
rect 41628 23238 41714 23290
rect 41766 23238 41852 23290
rect 41628 22954 41852 23238
rect 41628 22902 41714 22954
rect 41766 22902 41852 22954
rect 34136 22795 34192 22804
rect 34136 22730 34192 22739
rect 41628 22618 41852 22902
rect 41628 22566 41714 22618
rect 41766 22566 41852 22618
rect 41628 22284 41852 22566
rect 41628 22228 41712 22284
rect 41768 22228 41852 22284
rect 41628 21946 41852 22228
rect 41628 21894 41714 21946
rect 41766 21894 41852 21946
rect 41628 21610 41852 21894
rect 41628 21558 41714 21610
rect 41766 21558 41852 21610
rect 41628 21274 41852 21558
rect 41628 21222 41714 21274
rect 41766 21222 41852 21274
rect 41628 20938 41852 21222
rect 41628 20886 41714 20938
rect 41766 20886 41852 20938
rect 41628 20604 41852 20886
rect 41628 20548 41712 20604
rect 41768 20548 41852 20604
rect 41628 20266 41852 20548
rect 41628 20214 41714 20266
rect 41766 20214 41852 20266
rect 41628 19930 41852 20214
rect 41628 19878 41714 19930
rect 41766 19878 41852 19930
rect 41628 19594 41852 19878
rect 41628 19542 41714 19594
rect 41766 19542 41852 19594
rect 41628 19258 41852 19542
rect 41628 19206 41714 19258
rect 41766 19206 41852 19258
rect 41628 18924 41852 19206
rect 41628 18868 41712 18924
rect 41768 18868 41852 18924
rect 41628 18586 41852 18868
rect 41628 18534 41714 18586
rect 41766 18534 41852 18586
rect 41628 18250 41852 18534
rect 41628 18198 41714 18250
rect 41766 18198 41852 18250
rect 41628 17914 41852 18198
rect 41628 17862 41714 17914
rect 41766 17862 41852 17914
rect 41628 17578 41852 17862
rect 41628 17526 41714 17578
rect 41766 17526 41852 17578
rect 41628 17244 41852 17526
rect 41628 17188 41712 17244
rect 41768 17188 41852 17244
rect 41628 16906 41852 17188
rect 41628 16854 41714 16906
rect 41766 16854 41852 16906
rect 41628 16570 41852 16854
rect 41628 16518 41714 16570
rect 41766 16518 41852 16570
rect 41628 16234 41852 16518
rect 41628 16182 41714 16234
rect 41766 16182 41852 16234
rect 41628 15898 41852 16182
rect 41628 15846 41714 15898
rect 41766 15846 41852 15898
rect 41628 15564 41852 15846
rect 41628 15508 41712 15564
rect 41768 15508 41852 15564
rect 41628 15226 41852 15508
rect 41628 15174 41714 15226
rect 41766 15174 41852 15226
rect 41628 14890 41852 15174
rect 41628 14838 41714 14890
rect 41766 14838 41852 14890
rect 34052 14546 34108 14555
rect 15662 13242 15690 14527
rect 34052 14481 34108 14490
rect 41628 14554 41852 14838
rect 41628 14502 41714 14554
rect 41766 14502 41852 14554
rect 35134 14290 35190 14299
rect 33851 14219 33907 14228
rect 33851 14154 33907 14163
rect 34189 14219 34245 14228
rect 35134 14225 35190 14234
rect 34189 14154 34245 14163
rect 41628 14218 41852 14502
rect 41628 14166 41714 14218
rect 41766 14166 41852 14218
rect 41628 13884 41852 14166
rect 41628 13828 41712 13884
rect 41768 13828 41852 13884
rect 41628 13546 41852 13828
rect 41628 13494 41714 13546
rect 41766 13494 41852 13546
rect 15648 13233 15704 13242
rect 15648 13168 15704 13177
rect 41628 13210 41852 13494
rect 41628 13158 41714 13210
rect 41766 13158 41852 13210
rect 41628 12874 41852 13158
rect 40797 12859 40853 12868
rect 40797 12794 40853 12803
rect 41628 12822 41714 12874
rect 41766 12822 41852 12874
rect 33771 12661 33827 12670
rect 33771 12596 33827 12605
rect 34189 12661 34245 12670
rect 34189 12596 34245 12605
rect 35134 12590 35190 12599
rect 35134 12525 35190 12534
rect 41628 12538 41852 12822
rect 41628 12486 41714 12538
rect 41766 12486 41852 12538
rect 41628 12204 41852 12486
rect 41628 12148 41712 12204
rect 41768 12148 41852 12204
rect 41628 11866 41852 12148
rect 41628 11814 41714 11866
rect 41766 11814 41852 11866
rect 41628 11530 41852 11814
rect 41628 11478 41714 11530
rect 41766 11478 41852 11530
rect 35134 11462 35190 11471
rect 33691 11391 33747 11400
rect 33691 11326 33747 11335
rect 34189 11391 34245 11400
rect 35134 11397 35190 11406
rect 34189 11326 34245 11335
rect 41628 11194 41852 11478
rect 41628 11142 41714 11194
rect 41766 11142 41852 11194
rect 41628 10858 41852 11142
rect 41628 10806 41714 10858
rect 41766 10806 41852 10858
rect 19406 10677 19462 10686
rect 19406 10612 19462 10621
rect 20400 10677 20456 10686
rect 20400 10612 20456 10621
rect 20654 10677 20710 10686
rect 20654 10612 20710 10621
rect 21648 10677 21704 10686
rect 21648 10612 21704 10621
rect 21902 10677 21958 10686
rect 21902 10612 21958 10621
rect 22896 10677 22952 10686
rect 22896 10612 22952 10621
rect 23150 10677 23206 10686
rect 23150 10612 23206 10621
rect 24144 10677 24200 10686
rect 24144 10612 24200 10621
rect 41628 10524 41852 10806
rect 41628 10468 41712 10524
rect 41768 10468 41852 10524
rect 17299 10442 17355 10451
rect 17299 10377 17355 10386
rect 17313 6873 17341 10377
rect 41628 10186 41852 10468
rect 41628 10134 41714 10186
rect 41766 10134 41852 10186
rect 41628 9850 41852 10134
rect 33611 9833 33667 9842
rect 33611 9768 33667 9777
rect 34189 9833 34245 9842
rect 34189 9768 34245 9777
rect 41628 9798 41714 9850
rect 41766 9798 41852 9850
rect 35134 9762 35190 9771
rect 35134 9697 35190 9706
rect 41628 9514 41852 9798
rect 41628 9462 41714 9514
rect 41766 9462 41852 9514
rect 41628 9178 41852 9462
rect 41628 9126 41714 9178
rect 41766 9126 41852 9178
rect 17547 8991 17603 9000
rect 17547 8926 17603 8935
rect 17423 7593 17479 7602
rect 17423 7528 17479 7537
rect 17437 6873 17465 7528
rect 17561 6873 17589 8926
rect 41628 8844 41852 9126
rect 41628 8788 41712 8844
rect 41768 8788 41852 8844
rect 41628 8506 41852 8788
rect 41628 8454 41714 8506
rect 41766 8454 41852 8506
rect 41628 8170 41852 8454
rect 41628 8118 41714 8170
rect 41766 8118 41852 8170
rect 41628 7834 41852 8118
rect 41628 7782 41714 7834
rect 41766 7782 41852 7834
rect 41628 7498 41852 7782
rect 41628 7446 41714 7498
rect 41766 7446 41852 7498
rect 41628 7164 41852 7446
rect 41628 7108 41712 7164
rect 41768 7108 41852 7164
rect 9526 3307 9624 3321
rect 41628 6826 41852 7108
rect 41628 6774 41714 6826
rect 41766 6774 41852 6826
rect 41628 6490 41852 6774
rect 41628 6438 41714 6490
rect 41766 6438 41852 6490
rect 41628 6154 41852 6438
rect 41628 6102 41714 6154
rect 41766 6102 41852 6154
rect 41628 5818 41852 6102
rect 41628 5766 41714 5818
rect 41766 5766 41852 5818
rect 41628 5484 41852 5766
rect 41628 5428 41712 5484
rect 41768 5428 41852 5484
rect 41628 5146 41852 5428
rect 41628 5094 41714 5146
rect 41766 5094 41852 5146
rect 41628 4810 41852 5094
rect 41628 4758 41714 4810
rect 41766 4758 41852 4810
rect 41628 4474 41852 4758
rect 41628 4422 41714 4474
rect 41766 4422 41852 4474
rect 41628 4138 41852 4422
rect 41628 4086 41714 4138
rect 41766 4086 41852 4138
rect 41628 3804 41852 4086
rect 41628 3748 41712 3804
rect 41768 3748 41852 3804
rect 41628 3466 41852 3748
rect 41628 3414 41714 3466
rect 41766 3414 41852 3466
rect 6079 3297 6135 3306
rect 9526 3293 9647 3307
rect 6079 3232 6135 3241
rect 1646 3078 1732 3130
rect 1784 3078 1870 3130
rect 2858 3192 2914 3201
rect 2858 3127 2914 3136
rect 1646 2794 1870 3078
rect 9573 2936 9647 3293
rect 10836 3192 10892 3201
rect 10836 3127 10892 3136
rect 12004 3192 12060 3201
rect 12004 3127 12060 3136
rect 13172 3192 13228 3201
rect 13172 3127 13228 3136
rect 14340 3192 14396 3201
rect 14340 3127 14396 3136
rect 15508 3192 15564 3201
rect 15508 3127 15564 3136
rect 16676 3192 16732 3201
rect 16676 3127 16732 3136
rect 17844 3192 17900 3201
rect 17844 3127 17900 3136
rect 19012 3192 19068 3201
rect 19012 3127 19068 3136
rect 20180 3192 20236 3201
rect 20180 3127 20236 3136
rect 21348 3192 21404 3201
rect 21348 3127 21404 3136
rect 22516 3192 22572 3201
rect 22516 3127 22572 3136
rect 23684 3192 23740 3201
rect 23684 3127 23740 3136
rect 41628 3130 41852 3414
rect 9573 2908 9582 2936
rect 9638 2908 9647 2936
rect 41628 3078 41714 3130
rect 41766 3078 41852 3130
rect 9582 2871 9638 2880
rect 1646 2742 1732 2794
rect 1784 2742 1870 2794
rect 1646 2458 1870 2742
rect 1646 2406 1732 2458
rect 1784 2406 1870 2458
rect 1646 2124 1870 2406
rect 1646 2068 1730 2124
rect 1786 2068 1870 2124
rect 1646 1648 1870 2068
rect 41628 2794 41852 3078
rect 41628 2742 41714 2794
rect 41766 2742 41852 2794
rect 41628 2458 41852 2742
rect 41628 2406 41714 2458
rect 41766 2406 41852 2458
rect 41628 2124 41852 2406
rect 41628 2068 41712 2124
rect 41768 2068 41852 2124
rect 2066 1788 2122 1797
rect 2066 1723 2122 1732
rect 3746 1788 3802 1797
rect 3746 1723 3802 1732
rect 5426 1788 5482 1797
rect 5426 1723 5482 1732
rect 7106 1788 7162 1797
rect 7106 1723 7162 1732
rect 8786 1788 8842 1797
rect 8786 1723 8842 1732
rect 10466 1788 10522 1797
rect 10466 1723 10522 1732
rect 12146 1788 12202 1797
rect 12146 1723 12202 1732
rect 13826 1788 13882 1797
rect 13826 1723 13882 1732
rect 15506 1788 15562 1797
rect 15506 1723 15562 1732
rect 17186 1788 17242 1797
rect 17186 1723 17242 1732
rect 18866 1788 18922 1797
rect 18866 1723 18922 1732
rect 20546 1788 20602 1797
rect 20546 1723 20602 1732
rect 22226 1788 22282 1797
rect 22226 1723 22282 1732
rect 23906 1788 23962 1797
rect 23906 1723 23962 1732
rect 25586 1788 25642 1797
rect 25586 1723 25642 1732
rect 27266 1788 27322 1797
rect 27266 1723 27322 1732
rect 28946 1788 29002 1797
rect 28946 1723 29002 1732
rect 30626 1788 30682 1797
rect 30626 1723 30682 1732
rect 32306 1788 32362 1797
rect 32306 1723 32362 1732
rect 33986 1788 34042 1797
rect 33986 1723 34042 1732
rect 35666 1788 35722 1797
rect 35666 1723 35722 1732
rect 37346 1788 37402 1797
rect 37346 1723 37402 1732
rect 39026 1788 39082 1797
rect 39026 1723 39082 1732
rect 40706 1788 40762 1797
rect 40706 1723 40762 1732
rect 41628 1648 41852 2068
<< via2 >>
rect 2066 31410 2122 31412
rect 2066 31358 2068 31410
rect 2068 31358 2120 31410
rect 2120 31358 2122 31410
rect 2066 31356 2122 31358
rect 3746 31410 3802 31412
rect 3746 31358 3748 31410
rect 3748 31358 3800 31410
rect 3800 31358 3802 31410
rect 3746 31356 3802 31358
rect 5426 31410 5482 31412
rect 5426 31358 5428 31410
rect 5428 31358 5480 31410
rect 5480 31358 5482 31410
rect 5426 31356 5482 31358
rect 7106 31410 7162 31412
rect 7106 31358 7108 31410
rect 7108 31358 7160 31410
rect 7160 31358 7162 31410
rect 7106 31356 7162 31358
rect 8786 31410 8842 31412
rect 8786 31358 8788 31410
rect 8788 31358 8840 31410
rect 8840 31358 8842 31410
rect 8786 31356 8842 31358
rect 10466 31410 10522 31412
rect 10466 31358 10468 31410
rect 10468 31358 10520 31410
rect 10520 31358 10522 31410
rect 10466 31356 10522 31358
rect 12146 31410 12202 31412
rect 12146 31358 12148 31410
rect 12148 31358 12200 31410
rect 12200 31358 12202 31410
rect 12146 31356 12202 31358
rect 13826 31410 13882 31412
rect 13826 31358 13828 31410
rect 13828 31358 13880 31410
rect 13880 31358 13882 31410
rect 13826 31356 13882 31358
rect 15506 31410 15562 31412
rect 15506 31358 15508 31410
rect 15508 31358 15560 31410
rect 15560 31358 15562 31410
rect 15506 31356 15562 31358
rect 17186 31410 17242 31412
rect 17186 31358 17188 31410
rect 17188 31358 17240 31410
rect 17240 31358 17242 31410
rect 17186 31356 17242 31358
rect 18866 31410 18922 31412
rect 18866 31358 18868 31410
rect 18868 31358 18920 31410
rect 18920 31358 18922 31410
rect 18866 31356 18922 31358
rect 20546 31410 20602 31412
rect 20546 31358 20548 31410
rect 20548 31358 20600 31410
rect 20600 31358 20602 31410
rect 20546 31356 20602 31358
rect 22226 31410 22282 31412
rect 22226 31358 22228 31410
rect 22228 31358 22280 31410
rect 22280 31358 22282 31410
rect 22226 31356 22282 31358
rect 23906 31410 23962 31412
rect 23906 31358 23908 31410
rect 23908 31358 23960 31410
rect 23960 31358 23962 31410
rect 23906 31356 23962 31358
rect 25586 31410 25642 31412
rect 25586 31358 25588 31410
rect 25588 31358 25640 31410
rect 25640 31358 25642 31410
rect 25586 31356 25642 31358
rect 27266 31410 27322 31412
rect 27266 31358 27268 31410
rect 27268 31358 27320 31410
rect 27320 31358 27322 31410
rect 27266 31356 27322 31358
rect 28946 31410 29002 31412
rect 28946 31358 28948 31410
rect 28948 31358 29000 31410
rect 29000 31358 29002 31410
rect 28946 31356 29002 31358
rect 30626 31410 30682 31412
rect 30626 31358 30628 31410
rect 30628 31358 30680 31410
rect 30680 31358 30682 31410
rect 30626 31356 30682 31358
rect 32306 31410 32362 31412
rect 32306 31358 32308 31410
rect 32308 31358 32360 31410
rect 32360 31358 32362 31410
rect 32306 31356 32362 31358
rect 33986 31410 34042 31412
rect 33986 31358 33988 31410
rect 33988 31358 34040 31410
rect 34040 31358 34042 31410
rect 33986 31356 34042 31358
rect 35666 31410 35722 31412
rect 35666 31358 35668 31410
rect 35668 31358 35720 31410
rect 35720 31358 35722 31410
rect 35666 31356 35722 31358
rect 37346 31410 37402 31412
rect 37346 31358 37348 31410
rect 37348 31358 37400 31410
rect 37400 31358 37402 31410
rect 37346 31356 37402 31358
rect 39026 31410 39082 31412
rect 39026 31358 39028 31410
rect 39028 31358 39080 31410
rect 39080 31358 39082 31410
rect 39026 31356 39082 31358
rect 40706 31410 40762 31412
rect 40706 31358 40708 31410
rect 40708 31358 40760 31410
rect 40760 31358 40762 31410
rect 40706 31356 40762 31358
rect 1730 30682 1786 30684
rect 1730 30630 1732 30682
rect 1732 30630 1784 30682
rect 1784 30630 1786 30682
rect 1730 30628 1786 30630
rect 41712 30682 41768 30684
rect 41712 30630 41714 30682
rect 41714 30630 41766 30682
rect 41766 30630 41768 30682
rect 41712 30628 41768 30630
rect 40584 29952 40640 30008
rect 1730 29002 1786 29004
rect 1730 28950 1732 29002
rect 1732 28950 1784 29002
rect 1784 28950 1786 29002
rect 1730 28948 1786 28950
rect 1730 27322 1786 27324
rect 1730 27270 1732 27322
rect 1732 27270 1784 27322
rect 1784 27270 1786 27322
rect 1730 27268 1786 27270
rect 37447 29847 37503 29903
rect 8500 26206 8556 26262
rect 9445 26135 9501 26191
rect 9939 26189 9995 26191
rect 9939 26137 9941 26189
rect 9941 26137 9993 26189
rect 9993 26137 9995 26189
rect 9939 26135 9995 26137
rect 1730 25642 1786 25644
rect 1730 25590 1732 25642
rect 1732 25590 1784 25642
rect 1784 25590 1786 25642
rect 1730 25588 1786 25590
rect 25969 25551 26025 25607
rect 19406 25349 19462 25351
rect 19406 25297 19408 25349
rect 19408 25297 19460 25349
rect 19460 25297 19462 25349
rect 19406 25295 19462 25297
rect 20400 25349 20456 25351
rect 20400 25297 20402 25349
rect 20402 25297 20454 25349
rect 20454 25297 20456 25349
rect 20400 25295 20456 25297
rect 20654 25349 20710 25351
rect 20654 25297 20656 25349
rect 20656 25297 20708 25349
rect 20708 25297 20710 25349
rect 20654 25295 20710 25297
rect 21648 25349 21704 25351
rect 21648 25297 21650 25349
rect 21650 25297 21702 25349
rect 21702 25297 21704 25349
rect 21648 25295 21704 25297
rect 21902 25349 21958 25351
rect 21902 25297 21904 25349
rect 21904 25297 21956 25349
rect 21956 25297 21958 25349
rect 21902 25295 21958 25297
rect 22896 25349 22952 25351
rect 22896 25297 22898 25349
rect 22898 25297 22950 25349
rect 22950 25297 22952 25349
rect 22896 25295 22952 25297
rect 23150 25349 23206 25351
rect 23150 25297 23152 25349
rect 23152 25297 23204 25349
rect 23204 25297 23206 25349
rect 23150 25295 23206 25297
rect 24144 25349 24200 25351
rect 24144 25297 24146 25349
rect 24146 25297 24198 25349
rect 24198 25297 24200 25349
rect 24144 25295 24200 25297
rect 9445 24577 9501 24633
rect 9859 24631 9915 24633
rect 9859 24579 9861 24631
rect 9861 24579 9913 24631
rect 9913 24579 9915 24631
rect 9859 24577 9915 24579
rect 8500 24506 8556 24562
rect 26093 24190 26149 24246
rect 1730 23962 1786 23964
rect 1730 23910 1732 23962
rect 1732 23910 1784 23962
rect 1784 23910 1786 23962
rect 1730 23908 1786 23910
rect 8500 23378 8556 23434
rect 9445 23307 9501 23363
rect 9779 23361 9835 23363
rect 9779 23309 9781 23361
rect 9781 23309 9833 23361
rect 9833 23309 9835 23361
rect 9779 23307 9835 23309
rect 27902 22739 27958 22795
rect 1730 22282 1786 22284
rect 1730 22230 1732 22282
rect 1732 22230 1784 22282
rect 1784 22230 1786 22282
rect 1730 22228 1786 22230
rect 9445 21749 9501 21805
rect 9699 21803 9755 21805
rect 9699 21751 9701 21803
rect 9701 21751 9753 21803
rect 9753 21751 9755 21803
rect 9699 21749 9755 21751
rect 8500 21678 8556 21734
rect 9582 21422 9638 21478
rect 1730 20602 1786 20604
rect 1730 20550 1732 20602
rect 1732 20550 1784 20602
rect 1784 20550 1786 20602
rect 1730 20548 1786 20550
rect 2645 20285 2701 20341
rect 1730 18922 1786 18924
rect 1730 18870 1732 18922
rect 1732 18870 1784 18922
rect 1784 18870 1786 18922
rect 1730 18868 1786 18870
rect 1730 17242 1786 17244
rect 1730 17190 1732 17242
rect 1732 17190 1784 17242
rect 1784 17190 1786 17242
rect 1730 17188 1786 17190
rect 1730 15562 1786 15564
rect 1730 15510 1732 15562
rect 1732 15510 1784 15562
rect 1784 15510 1786 15562
rect 1730 15508 1786 15510
rect 1730 13882 1786 13884
rect 1730 13830 1732 13882
rect 1732 13830 1784 13882
rect 1784 13830 1786 13882
rect 1730 13828 1786 13830
rect 9498 13177 9554 13233
rect 1730 12202 1786 12204
rect 1730 12150 1732 12202
rect 1732 12150 1784 12202
rect 1784 12150 1786 12202
rect 1730 12148 1786 12150
rect 1730 10522 1786 10524
rect 1730 10470 1732 10522
rect 1732 10470 1784 10522
rect 1784 10470 1786 10522
rect 1730 10468 1786 10470
rect 9498 10386 9554 10442
rect 9498 8935 9554 8991
rect 1730 8842 1786 8844
rect 1730 8790 1732 8842
rect 1732 8790 1784 8842
rect 1784 8790 1786 8842
rect 1730 8788 1786 8790
rect 9498 7537 9554 7593
rect 1730 7162 1786 7164
rect 1730 7110 1732 7162
rect 1732 7110 1784 7162
rect 1784 7110 1786 7162
rect 1730 7108 1786 7110
rect 1730 5482 1786 5484
rect 1730 5430 1732 5482
rect 1732 5430 1784 5482
rect 1784 5430 1786 5482
rect 1730 5428 1786 5430
rect 2858 4836 2914 4892
rect 1730 3802 1786 3804
rect 1730 3750 1732 3802
rect 1732 3750 1784 3802
rect 1784 3750 1786 3802
rect 1730 3748 1786 3750
rect 41712 29002 41768 29004
rect 41712 28950 41714 29002
rect 41714 28950 41766 29002
rect 41766 28950 41768 29002
rect 41712 28948 41768 28950
rect 41712 27322 41768 27324
rect 41712 27270 41714 27322
rect 41714 27270 41766 27322
rect 41766 27270 41768 27322
rect 41712 27268 41768 27270
rect 34136 25551 34192 25607
rect 41712 25642 41768 25644
rect 41712 25590 41714 25642
rect 41714 25590 41766 25642
rect 41766 25590 41768 25642
rect 41712 25588 41768 25590
rect 34136 24190 34192 24246
rect 41712 23962 41768 23964
rect 41712 23910 41714 23962
rect 41714 23910 41766 23962
rect 41766 23910 41768 23962
rect 41712 23908 41768 23910
rect 34136 22739 34192 22795
rect 41712 22282 41768 22284
rect 41712 22230 41714 22282
rect 41714 22230 41766 22282
rect 41766 22230 41768 22282
rect 41712 22228 41768 22230
rect 41712 20602 41768 20604
rect 41712 20550 41714 20602
rect 41714 20550 41766 20602
rect 41766 20550 41768 20602
rect 41712 20548 41768 20550
rect 41712 18922 41768 18924
rect 41712 18870 41714 18922
rect 41714 18870 41766 18922
rect 41766 18870 41768 18922
rect 41712 18868 41768 18870
rect 41712 17242 41768 17244
rect 41712 17190 41714 17242
rect 41714 17190 41766 17242
rect 41766 17190 41768 17242
rect 41712 17188 41768 17190
rect 41712 15562 41768 15564
rect 41712 15510 41714 15562
rect 41714 15510 41766 15562
rect 41766 15510 41768 15562
rect 41712 15508 41768 15510
rect 34052 14490 34108 14546
rect 35134 14234 35190 14290
rect 33851 14217 33907 14219
rect 33851 14165 33853 14217
rect 33853 14165 33905 14217
rect 33905 14165 33907 14217
rect 33851 14163 33907 14165
rect 34189 14163 34245 14219
rect 41712 13882 41768 13884
rect 41712 13830 41714 13882
rect 41714 13830 41766 13882
rect 41766 13830 41768 13882
rect 41712 13828 41768 13830
rect 15648 13177 15704 13233
rect 40797 12803 40853 12859
rect 33771 12659 33827 12661
rect 33771 12607 33773 12659
rect 33773 12607 33825 12659
rect 33825 12607 33827 12659
rect 33771 12605 33827 12607
rect 34189 12605 34245 12661
rect 35134 12534 35190 12590
rect 41712 12202 41768 12204
rect 41712 12150 41714 12202
rect 41714 12150 41766 12202
rect 41766 12150 41768 12202
rect 41712 12148 41768 12150
rect 35134 11406 35190 11462
rect 33691 11389 33747 11391
rect 33691 11337 33693 11389
rect 33693 11337 33745 11389
rect 33745 11337 33747 11389
rect 33691 11335 33747 11337
rect 34189 11335 34245 11391
rect 19406 10675 19462 10677
rect 19406 10623 19408 10675
rect 19408 10623 19460 10675
rect 19460 10623 19462 10675
rect 19406 10621 19462 10623
rect 20400 10675 20456 10677
rect 20400 10623 20402 10675
rect 20402 10623 20454 10675
rect 20454 10623 20456 10675
rect 20400 10621 20456 10623
rect 20654 10675 20710 10677
rect 20654 10623 20656 10675
rect 20656 10623 20708 10675
rect 20708 10623 20710 10675
rect 20654 10621 20710 10623
rect 21648 10675 21704 10677
rect 21648 10623 21650 10675
rect 21650 10623 21702 10675
rect 21702 10623 21704 10675
rect 21648 10621 21704 10623
rect 21902 10675 21958 10677
rect 21902 10623 21904 10675
rect 21904 10623 21956 10675
rect 21956 10623 21958 10675
rect 21902 10621 21958 10623
rect 22896 10675 22952 10677
rect 22896 10623 22898 10675
rect 22898 10623 22950 10675
rect 22950 10623 22952 10675
rect 22896 10621 22952 10623
rect 23150 10675 23206 10677
rect 23150 10623 23152 10675
rect 23152 10623 23204 10675
rect 23204 10623 23206 10675
rect 23150 10621 23206 10623
rect 24144 10675 24200 10677
rect 24144 10623 24146 10675
rect 24146 10623 24198 10675
rect 24198 10623 24200 10675
rect 24144 10621 24200 10623
rect 41712 10522 41768 10524
rect 41712 10470 41714 10522
rect 41714 10470 41766 10522
rect 41766 10470 41768 10522
rect 41712 10468 41768 10470
rect 17299 10386 17355 10442
rect 33611 9831 33667 9833
rect 33611 9779 33613 9831
rect 33613 9779 33665 9831
rect 33665 9779 33667 9831
rect 33611 9777 33667 9779
rect 34189 9777 34245 9833
rect 35134 9706 35190 9762
rect 17547 8935 17603 8991
rect 17423 7537 17479 7593
rect 41712 8842 41768 8844
rect 41712 8790 41714 8842
rect 41714 8790 41766 8842
rect 41766 8790 41768 8842
rect 41712 8788 41768 8790
rect 41712 7162 41768 7164
rect 41712 7110 41714 7162
rect 41714 7110 41766 7162
rect 41766 7110 41768 7162
rect 41712 7108 41768 7110
rect 41712 5482 41768 5484
rect 41712 5430 41714 5482
rect 41714 5430 41766 5482
rect 41766 5430 41768 5482
rect 41712 5428 41768 5430
rect 41712 3802 41768 3804
rect 41712 3750 41714 3802
rect 41714 3750 41766 3802
rect 41766 3750 41768 3802
rect 41712 3748 41768 3750
rect 6079 3241 6135 3297
rect 2858 3136 2914 3192
rect 10836 3136 10892 3192
rect 12004 3136 12060 3192
rect 13172 3136 13228 3192
rect 14340 3136 14396 3192
rect 15508 3136 15564 3192
rect 16676 3136 16732 3192
rect 17844 3136 17900 3192
rect 19012 3136 19068 3192
rect 20180 3136 20236 3192
rect 21348 3136 21404 3192
rect 22516 3136 22572 3192
rect 23684 3136 23740 3192
rect 9582 2880 9638 2936
rect 1730 2122 1786 2124
rect 1730 2070 1732 2122
rect 1732 2070 1784 2122
rect 1784 2070 1786 2122
rect 1730 2068 1786 2070
rect 41712 2122 41768 2124
rect 41712 2070 41714 2122
rect 41714 2070 41766 2122
rect 41766 2070 41768 2122
rect 41712 2068 41768 2070
rect 2066 1786 2122 1788
rect 2066 1734 2068 1786
rect 2068 1734 2120 1786
rect 2120 1734 2122 1786
rect 2066 1732 2122 1734
rect 3746 1786 3802 1788
rect 3746 1734 3748 1786
rect 3748 1734 3800 1786
rect 3800 1734 3802 1786
rect 3746 1732 3802 1734
rect 5426 1786 5482 1788
rect 5426 1734 5428 1786
rect 5428 1734 5480 1786
rect 5480 1734 5482 1786
rect 5426 1732 5482 1734
rect 7106 1786 7162 1788
rect 7106 1734 7108 1786
rect 7108 1734 7160 1786
rect 7160 1734 7162 1786
rect 7106 1732 7162 1734
rect 8786 1786 8842 1788
rect 8786 1734 8788 1786
rect 8788 1734 8840 1786
rect 8840 1734 8842 1786
rect 8786 1732 8842 1734
rect 10466 1786 10522 1788
rect 10466 1734 10468 1786
rect 10468 1734 10520 1786
rect 10520 1734 10522 1786
rect 10466 1732 10522 1734
rect 12146 1786 12202 1788
rect 12146 1734 12148 1786
rect 12148 1734 12200 1786
rect 12200 1734 12202 1786
rect 12146 1732 12202 1734
rect 13826 1786 13882 1788
rect 13826 1734 13828 1786
rect 13828 1734 13880 1786
rect 13880 1734 13882 1786
rect 13826 1732 13882 1734
rect 15506 1786 15562 1788
rect 15506 1734 15508 1786
rect 15508 1734 15560 1786
rect 15560 1734 15562 1786
rect 15506 1732 15562 1734
rect 17186 1786 17242 1788
rect 17186 1734 17188 1786
rect 17188 1734 17240 1786
rect 17240 1734 17242 1786
rect 17186 1732 17242 1734
rect 18866 1786 18922 1788
rect 18866 1734 18868 1786
rect 18868 1734 18920 1786
rect 18920 1734 18922 1786
rect 18866 1732 18922 1734
rect 20546 1786 20602 1788
rect 20546 1734 20548 1786
rect 20548 1734 20600 1786
rect 20600 1734 20602 1786
rect 20546 1732 20602 1734
rect 22226 1786 22282 1788
rect 22226 1734 22228 1786
rect 22228 1734 22280 1786
rect 22280 1734 22282 1786
rect 22226 1732 22282 1734
rect 23906 1786 23962 1788
rect 23906 1734 23908 1786
rect 23908 1734 23960 1786
rect 23960 1734 23962 1786
rect 23906 1732 23962 1734
rect 25586 1786 25642 1788
rect 25586 1734 25588 1786
rect 25588 1734 25640 1786
rect 25640 1734 25642 1786
rect 25586 1732 25642 1734
rect 27266 1786 27322 1788
rect 27266 1734 27268 1786
rect 27268 1734 27320 1786
rect 27320 1734 27322 1786
rect 27266 1732 27322 1734
rect 28946 1786 29002 1788
rect 28946 1734 28948 1786
rect 28948 1734 29000 1786
rect 29000 1734 29002 1786
rect 28946 1732 29002 1734
rect 30626 1786 30682 1788
rect 30626 1734 30628 1786
rect 30628 1734 30680 1786
rect 30680 1734 30682 1786
rect 30626 1732 30682 1734
rect 32306 1786 32362 1788
rect 32306 1734 32308 1786
rect 32308 1734 32360 1786
rect 32360 1734 32362 1786
rect 32306 1732 32362 1734
rect 33986 1786 34042 1788
rect 33986 1734 33988 1786
rect 33988 1734 34040 1786
rect 34040 1734 34042 1786
rect 33986 1732 34042 1734
rect 35666 1786 35722 1788
rect 35666 1734 35668 1786
rect 35668 1734 35720 1786
rect 35720 1734 35722 1786
rect 35666 1732 35722 1734
rect 37346 1786 37402 1788
rect 37346 1734 37348 1786
rect 37348 1734 37400 1786
rect 37400 1734 37402 1786
rect 37346 1732 37402 1734
rect 39026 1786 39082 1788
rect 39026 1734 39028 1786
rect 39028 1734 39080 1786
rect 39080 1734 39082 1786
rect 39026 1732 39082 1734
rect 40706 1786 40762 1788
rect 40706 1734 40708 1786
rect 40708 1734 40760 1786
rect 40760 1734 40762 1786
rect 40706 1732 40762 1734
<< metal3 >>
rect 272 32846 43188 32852
rect 272 32782 278 32846
rect 342 32782 414 32846
rect 478 32782 550 32846
rect 614 32782 42846 32846
rect 42910 32782 42982 32846
rect 43046 32782 43118 32846
rect 43182 32782 43188 32846
rect 272 32710 43188 32782
rect 272 32646 278 32710
rect 342 32646 414 32710
rect 478 32646 550 32710
rect 614 32646 42846 32710
rect 42910 32646 42982 32710
rect 43046 32646 43118 32710
rect 43182 32646 43188 32710
rect 272 32574 43188 32646
rect 272 32510 278 32574
rect 342 32510 414 32574
rect 478 32510 550 32574
rect 614 32510 34278 32574
rect 34342 32510 42846 32574
rect 42910 32510 42982 32574
rect 43046 32510 43118 32574
rect 43182 32510 43188 32574
rect 272 32504 43188 32510
rect 952 32166 42508 32172
rect 952 32102 958 32166
rect 1022 32102 1094 32166
rect 1158 32102 1230 32166
rect 1294 32102 42166 32166
rect 42230 32102 42302 32166
rect 42366 32102 42438 32166
rect 42502 32102 42508 32166
rect 952 32030 42508 32102
rect 952 31966 958 32030
rect 1022 31966 1094 32030
rect 1158 31966 1230 32030
rect 1294 31966 42166 32030
rect 42230 31966 42302 32030
rect 42366 31966 42438 32030
rect 42502 31966 42508 32030
rect 952 31894 42508 31966
rect 952 31830 958 31894
rect 1022 31830 1094 31894
rect 1158 31830 1230 31894
rect 1294 31830 2182 31894
rect 2246 31830 3814 31894
rect 3878 31830 5310 31894
rect 5374 31830 7078 31894
rect 7142 31830 8710 31894
rect 8774 31830 10342 31894
rect 10406 31830 12110 31894
rect 12174 31830 13742 31894
rect 13806 31830 15646 31894
rect 15710 31830 17278 31894
rect 17342 31830 18774 31894
rect 18838 31830 20270 31894
rect 20334 31830 22310 31894
rect 22374 31830 23806 31894
rect 23870 31830 25574 31894
rect 25638 31830 27206 31894
rect 27270 31830 28974 31894
rect 29038 31830 30606 31894
rect 30670 31830 32238 31894
rect 32302 31830 34006 31894
rect 34070 31830 35638 31894
rect 35702 31830 37270 31894
rect 37334 31830 38902 31894
rect 38966 31830 40670 31894
rect 40734 31830 42166 31894
rect 42230 31830 42302 31894
rect 42366 31830 42438 31894
rect 42502 31830 42508 31894
rect 952 31824 42508 31830
rect 2040 31486 2252 31492
rect 2040 31422 2182 31486
rect 2246 31422 2252 31486
rect 2040 31412 2252 31422
rect 2040 31356 2066 31412
rect 2122 31356 2252 31412
rect 2040 31280 2252 31356
rect 3672 31486 3884 31492
rect 3672 31422 3814 31486
rect 3878 31422 3884 31486
rect 3672 31412 3884 31422
rect 3672 31356 3746 31412
rect 3802 31356 3884 31412
rect 3672 31280 3884 31356
rect 5304 31486 5516 31492
rect 5304 31422 5310 31486
rect 5374 31422 5516 31486
rect 5304 31412 5516 31422
rect 5304 31356 5426 31412
rect 5482 31356 5516 31412
rect 5304 31280 5516 31356
rect 7072 31486 7284 31492
rect 7072 31422 7078 31486
rect 7142 31422 7284 31486
rect 7072 31412 7284 31422
rect 7072 31356 7106 31412
rect 7162 31356 7284 31412
rect 7072 31280 7284 31356
rect 8704 31486 8916 31492
rect 8704 31422 8710 31486
rect 8774 31422 8916 31486
rect 8704 31412 8916 31422
rect 8704 31356 8786 31412
rect 8842 31356 8916 31412
rect 8704 31280 8916 31356
rect 10336 31486 10548 31492
rect 10336 31422 10342 31486
rect 10406 31422 10548 31486
rect 10336 31412 10548 31422
rect 10336 31356 10466 31412
rect 10522 31356 10548 31412
rect 10336 31280 10548 31356
rect 12104 31486 12316 31492
rect 12104 31422 12110 31486
rect 12174 31422 12316 31486
rect 12104 31412 12316 31422
rect 12104 31356 12146 31412
rect 12202 31356 12316 31412
rect 12104 31280 12316 31356
rect 13736 31486 13948 31492
rect 13736 31422 13742 31486
rect 13806 31422 13948 31486
rect 13736 31412 13948 31422
rect 13736 31356 13826 31412
rect 13882 31356 13948 31412
rect 13736 31280 13948 31356
rect 15368 31486 15716 31492
rect 15368 31422 15646 31486
rect 15710 31422 15716 31486
rect 15368 31412 15716 31422
rect 15368 31356 15506 31412
rect 15562 31356 15716 31412
rect 15368 31280 15716 31356
rect 17136 31486 17348 31492
rect 17136 31422 17278 31486
rect 17342 31422 17348 31486
rect 17136 31412 17348 31422
rect 17136 31356 17186 31412
rect 17242 31356 17348 31412
rect 17136 31280 17348 31356
rect 18768 31486 18980 31492
rect 18768 31422 18774 31486
rect 18838 31422 18980 31486
rect 18768 31412 18980 31422
rect 20264 31486 20748 31492
rect 20264 31422 20270 31486
rect 20334 31422 20748 31486
rect 20264 31416 20748 31422
rect 18768 31356 18866 31412
rect 18922 31356 18980 31412
rect 18768 31280 18980 31356
rect 20400 31412 20748 31416
rect 20400 31356 20546 31412
rect 20602 31356 20748 31412
rect 20400 31280 20748 31356
rect 22168 31486 22380 31492
rect 22168 31422 22310 31486
rect 22374 31422 22380 31486
rect 22168 31412 22380 31422
rect 22168 31356 22226 31412
rect 22282 31356 22380 31412
rect 22168 31280 22380 31356
rect 23800 31486 24012 31492
rect 23800 31422 23806 31486
rect 23870 31422 24012 31486
rect 23800 31412 24012 31422
rect 23800 31356 23906 31412
rect 23962 31356 24012 31412
rect 23800 31280 24012 31356
rect 25432 31486 25780 31492
rect 25432 31422 25574 31486
rect 25638 31422 25780 31486
rect 25432 31412 25780 31422
rect 25432 31356 25586 31412
rect 25642 31356 25780 31412
rect 25432 31280 25780 31356
rect 27200 31486 27412 31492
rect 27200 31422 27206 31486
rect 27270 31422 27412 31486
rect 27200 31412 27412 31422
rect 27200 31356 27266 31412
rect 27322 31356 27412 31412
rect 27200 31280 27412 31356
rect 28832 31486 29044 31492
rect 28832 31422 28974 31486
rect 29038 31422 29044 31486
rect 28832 31412 29044 31422
rect 28832 31356 28946 31412
rect 29002 31356 29044 31412
rect 28832 31280 29044 31356
rect 30600 31486 30812 31492
rect 30600 31422 30606 31486
rect 30670 31422 30812 31486
rect 30600 31412 30812 31422
rect 30600 31356 30626 31412
rect 30682 31356 30812 31412
rect 30600 31280 30812 31356
rect 32232 31486 32444 31492
rect 32232 31422 32238 31486
rect 32302 31422 32444 31486
rect 32232 31412 32444 31422
rect 32232 31356 32306 31412
rect 32362 31356 32444 31412
rect 32232 31280 32444 31356
rect 33864 31486 34076 31492
rect 33864 31422 34006 31486
rect 34070 31422 34076 31486
rect 33864 31412 34076 31422
rect 33864 31356 33986 31412
rect 34042 31356 34076 31412
rect 35632 31486 35844 31492
rect 35632 31422 35638 31486
rect 35702 31422 35844 31486
rect 35632 31412 35844 31422
rect 35632 31356 35666 31412
rect 35722 31356 35844 31412
rect 33864 31350 34212 31356
rect 33864 31286 34142 31350
rect 34206 31286 34212 31350
rect 33864 31280 34212 31286
rect 35632 31280 35844 31356
rect 37264 31486 37476 31492
rect 37264 31422 37270 31486
rect 37334 31422 37476 31486
rect 37264 31412 37476 31422
rect 37264 31356 37346 31412
rect 37402 31356 37476 31412
rect 37264 31280 37476 31356
rect 38896 31486 39108 31492
rect 38896 31422 38902 31486
rect 38966 31422 39108 31486
rect 38896 31412 39108 31422
rect 38896 31356 39026 31412
rect 39082 31356 39108 31412
rect 38896 31280 39108 31356
rect 40664 31486 40876 31492
rect 40664 31422 40670 31486
rect 40734 31422 40876 31486
rect 40664 31412 40876 31422
rect 40664 31356 40706 31412
rect 40762 31356 40876 31412
rect 40664 31280 40876 31356
rect 1224 30806 1844 30812
rect 1224 30742 1230 30806
rect 1294 30742 1844 30806
rect 1224 30736 1844 30742
rect 1632 30684 1844 30736
rect 1632 30628 1730 30684
rect 1786 30628 1844 30684
rect 41616 30806 42236 30812
rect 41616 30742 42166 30806
rect 42230 30742 42236 30806
rect 41616 30736 42236 30742
rect 41616 30684 41828 30736
rect 1632 30600 1844 30628
rect 34136 30670 34348 30676
rect 34136 30606 34278 30670
rect 34342 30606 34348 30670
rect 34136 30540 34348 30606
rect 34000 30534 34348 30540
rect 34000 30470 34006 30534
rect 34070 30470 34348 30534
rect 34000 30464 34348 30470
rect 40664 30540 40876 30676
rect 41616 30628 41712 30684
rect 41768 30628 41828 30684
rect 41616 30600 41828 30628
rect 40664 30534 42916 30540
rect 40664 30470 42846 30534
rect 42910 30470 42916 30534
rect 40664 30464 42916 30470
rect 40528 30056 43460 30132
rect 40528 30008 40740 30056
rect 37400 29990 37612 29996
rect 37400 29926 37406 29990
rect 37470 29926 37612 29990
rect 37400 29903 37612 29926
rect 40528 29952 40584 30008
rect 40640 29952 40740 30008
rect 40528 29920 40740 29952
rect 37400 29847 37447 29903
rect 37503 29847 37612 29903
rect 37400 29784 37612 29847
rect 34136 29174 34348 29180
rect 34136 29110 34142 29174
rect 34206 29110 34348 29174
rect 1632 29004 1844 29044
rect 1632 28948 1730 29004
rect 1786 28948 1844 29004
rect 34136 29038 34348 29110
rect 34136 28974 34278 29038
rect 34342 28974 34348 29038
rect 34136 28968 34348 28974
rect 40664 29044 40876 29180
rect 40664 29004 41828 29044
rect 40664 28968 41712 29004
rect 1632 28908 1844 28948
rect 1224 28902 1844 28908
rect 1224 28838 1230 28902
rect 1294 28838 1844 28902
rect 1224 28832 1844 28838
rect 41616 28948 41712 28968
rect 41768 28948 41828 29004
rect 41616 28908 41828 28948
rect 41616 28902 42236 28908
rect 41616 28838 42166 28902
rect 42230 28838 42236 28902
rect 41616 28832 42236 28838
rect 34038 27814 34348 27820
rect 34000 27750 34006 27814
rect 34070 27750 34348 27814
rect 34038 27744 34348 27750
rect 34136 27684 34348 27744
rect 34136 27678 34446 27684
rect 34136 27614 34414 27678
rect 34478 27614 34484 27678
rect 34136 27608 34446 27614
rect 1224 27406 1844 27412
rect 1224 27342 1230 27406
rect 1294 27342 1844 27406
rect 1224 27336 1844 27342
rect 1632 27324 1844 27336
rect 1632 27268 1730 27324
rect 1786 27268 1844 27324
rect 1632 27200 1844 27268
rect 41616 27406 42236 27412
rect 41616 27342 42166 27406
rect 42230 27342 42236 27406
rect 41616 27336 42236 27342
rect 41616 27324 41828 27336
rect 41616 27268 41712 27324
rect 41768 27268 41828 27324
rect 41616 27200 41828 27268
rect 8840 26726 9052 26868
rect 8840 26662 8846 26726
rect 8910 26662 9052 26726
rect 8840 26656 9052 26662
rect 34136 26454 34348 26460
rect 34136 26390 34278 26454
rect 34342 26390 34348 26454
rect 8432 26318 8644 26324
rect 8432 26262 8574 26318
rect 8432 26206 8500 26262
rect 8556 26254 8574 26262
rect 8638 26254 8644 26318
rect 8556 26206 8644 26254
rect 34136 26318 34348 26390
rect 34136 26254 34142 26318
rect 34206 26254 34348 26318
rect 34136 26248 34348 26254
rect 8432 26112 8644 26206
rect 9440 26193 9506 26196
rect 9934 26193 10000 26196
rect 9440 26191 10000 26193
rect 9440 26135 9445 26191
rect 9501 26135 9939 26191
rect 9995 26135 10000 26191
rect 9440 26133 10000 26135
rect 9440 26130 9506 26133
rect 9934 26130 10000 26133
rect 1632 25644 1844 25780
rect 20166 25774 21020 25780
rect 21526 25774 22244 25780
rect 22750 25774 23468 25780
rect 20128 25710 20134 25774
rect 20198 25710 20950 25774
rect 21014 25710 21020 25774
rect 21488 25710 21494 25774
rect 21558 25710 22174 25774
rect 22238 25710 22244 25774
rect 22712 25710 22718 25774
rect 22782 25710 23398 25774
rect 23462 25710 23468 25774
rect 20166 25704 21020 25710
rect 21526 25704 22244 25710
rect 22750 25704 23468 25710
rect 1224 25638 1730 25644
rect 1224 25574 1230 25638
rect 1294 25588 1730 25638
rect 1786 25588 1844 25644
rect 41616 25644 41828 25780
rect 1294 25574 1844 25588
rect 1224 25568 1844 25574
rect 1632 25432 1844 25568
rect 25964 25609 26030 25612
rect 34131 25609 34197 25612
rect 25964 25607 34197 25609
rect 25964 25551 25969 25607
rect 26025 25551 34136 25607
rect 34192 25551 34197 25607
rect 25964 25549 34197 25551
rect 25964 25546 26030 25549
rect 34131 25546 34197 25549
rect 41616 25588 41712 25644
rect 41768 25588 41828 25644
rect 41616 25508 41828 25588
rect 8840 25366 9052 25508
rect 8840 25302 8982 25366
rect 9046 25302 9052 25366
rect 8840 25296 9052 25302
rect 19312 25502 19524 25508
rect 19312 25438 19318 25502
rect 19382 25438 19524 25502
rect 19312 25351 19524 25438
rect 19720 25391 19796 25508
rect 19312 25295 19406 25351
rect 19462 25295 19524 25351
rect 19312 25160 19524 25295
rect 19639 25372 19796 25391
rect 19992 25502 20204 25508
rect 19992 25438 20134 25502
rect 20198 25438 20204 25502
rect 19992 25391 20204 25438
rect 20400 25502 20476 25508
rect 20400 25438 20406 25502
rect 20470 25438 20476 25502
rect 19992 25372 20223 25391
rect 20400 25372 20476 25438
rect 20672 25502 20748 25508
rect 20672 25438 20678 25502
rect 20742 25438 20748 25502
rect 20672 25372 20748 25438
rect 20944 25502 21020 25508
rect 20944 25438 20950 25502
rect 21014 25438 21020 25502
rect 20944 25391 21020 25438
rect 19639 25296 20223 25372
rect 19639 25293 19796 25296
rect 19720 25160 19796 25293
rect 19992 25293 20223 25296
rect 20379 25351 20477 25372
rect 20379 25295 20400 25351
rect 20456 25295 20477 25351
rect 20536 25351 20748 25372
rect 20536 25296 20654 25351
rect 19992 25160 20204 25293
rect 20379 25274 20477 25295
rect 20633 25295 20654 25296
rect 20710 25295 20748 25351
rect 20633 25274 20748 25295
rect 20887 25293 21020 25391
rect 20400 25160 20476 25274
rect 20672 25160 20748 25274
rect 20944 25236 21020 25293
rect 21352 25502 21564 25508
rect 21352 25438 21494 25502
rect 21558 25438 21564 25502
rect 21352 25236 21564 25438
rect 20944 25160 21564 25236
rect 21624 25502 21700 25508
rect 21624 25438 21630 25502
rect 21694 25438 21700 25502
rect 21624 25372 21700 25438
rect 21896 25502 21972 25508
rect 21896 25438 21902 25502
rect 21966 25438 21972 25502
rect 21896 25372 21972 25438
rect 22168 25502 22788 25508
rect 22168 25438 22174 25502
rect 22238 25438 22718 25502
rect 22782 25438 22788 25502
rect 22168 25432 22788 25438
rect 22168 25391 22244 25432
rect 21624 25351 21725 25372
rect 21624 25295 21648 25351
rect 21704 25295 21725 25351
rect 21624 25274 21725 25295
rect 21881 25351 21979 25372
rect 21881 25295 21902 25351
rect 21958 25295 21979 25351
rect 21881 25274 21979 25295
rect 22135 25293 22244 25391
rect 21624 25160 21700 25274
rect 21896 25160 21972 25274
rect 22168 25160 22244 25293
rect 22576 25160 22788 25432
rect 22848 25502 23060 25508
rect 22848 25438 22854 25502
rect 22918 25438 23060 25502
rect 22848 25351 23060 25438
rect 22848 25295 22896 25351
rect 22952 25295 23060 25351
rect 22848 25160 23060 25295
rect 23120 25502 23196 25508
rect 23120 25438 23126 25502
rect 23190 25438 23196 25502
rect 23120 25372 23196 25438
rect 23392 25502 23604 25508
rect 23392 25438 23398 25502
rect 23462 25438 23604 25502
rect 23392 25391 23604 25438
rect 23383 25372 23604 25391
rect 23800 25372 24012 25508
rect 23120 25351 23227 25372
rect 23120 25295 23150 25351
rect 23206 25295 23227 25351
rect 23120 25274 23227 25295
rect 23383 25296 24012 25372
rect 23383 25293 23604 25296
rect 23120 25160 23196 25274
rect 23392 25160 23604 25293
rect 23800 25230 24012 25296
rect 23800 25166 23942 25230
rect 24006 25166 24012 25230
rect 23800 25160 24012 25166
rect 24072 25502 24284 25508
rect 24072 25438 24214 25502
rect 24278 25438 24284 25502
rect 24072 25351 24284 25438
rect 41616 25502 42236 25508
rect 41616 25438 42166 25502
rect 42230 25438 42236 25502
rect 41616 25432 42236 25438
rect 24072 25295 24144 25351
rect 24200 25295 24284 25351
rect 24072 25160 24284 25295
rect 19584 25024 20340 25100
rect 19584 24888 19796 25024
rect 19992 24964 20340 25024
rect 20808 24964 21020 25100
rect 21352 24964 21564 25100
rect 22032 25024 24012 25100
rect 22032 24964 22244 25024
rect 19992 24958 22244 24964
rect 19992 24894 21494 24958
rect 21558 24894 22244 24958
rect 19992 24888 22244 24894
rect 22576 24958 22788 25024
rect 22576 24894 22582 24958
rect 22646 24894 22788 24958
rect 22576 24888 22788 24894
rect 23256 24888 23604 25024
rect 23800 24888 24012 25024
rect 34136 24958 34484 24964
rect 34136 24894 34414 24958
rect 34478 24894 34484 24958
rect 34136 24888 34484 24894
rect 39304 24888 40196 24964
rect 34136 24822 34348 24888
rect 34136 24758 34278 24822
rect 34342 24758 34348 24822
rect 34136 24752 34348 24758
rect 39304 24752 39516 24888
rect 39984 24828 40196 24888
rect 39984 24822 41692 24828
rect 39984 24758 41622 24822
rect 41686 24758 41692 24822
rect 39984 24752 41692 24758
rect 0 24616 8644 24692
rect 8432 24562 8644 24616
rect 9440 24635 9506 24638
rect 9854 24635 9920 24638
rect 9440 24633 9920 24635
rect 9440 24577 9445 24633
rect 9501 24577 9859 24633
rect 9915 24577 9920 24633
rect 9440 24575 9920 24577
rect 9440 24572 9506 24575
rect 9854 24572 9920 24575
rect 8432 24506 8500 24562
rect 8556 24506 8644 24562
rect 8432 24480 8644 24506
rect 19584 24208 20340 24284
rect 8840 24142 9052 24148
rect 8840 24078 8846 24142
rect 8910 24078 9052 24142
rect 1632 23964 1844 24012
rect 1632 23908 1730 23964
rect 1786 23908 1844 23964
rect 1632 23876 1844 23908
rect 1224 23870 1844 23876
rect 1224 23806 1230 23870
rect 1294 23806 1844 23870
rect 1224 23800 1844 23806
rect 8840 23870 9052 24078
rect 19584 24142 19796 24208
rect 19584 24078 19590 24142
rect 19654 24078 19796 24142
rect 19584 24072 19796 24078
rect 20128 24148 20340 24208
rect 20808 24148 21020 24284
rect 21352 24278 21564 24284
rect 21352 24214 21494 24278
rect 21558 24214 21564 24278
rect 21352 24148 21564 24214
rect 20128 24072 21564 24148
rect 22032 24148 22244 24284
rect 22576 24278 23604 24284
rect 22576 24214 22582 24278
rect 22646 24214 23604 24278
rect 22576 24208 23604 24214
rect 22576 24148 22788 24208
rect 22032 24072 22788 24148
rect 23256 24148 23604 24208
rect 23800 24148 24012 24284
rect 26088 24248 26154 24251
rect 34131 24248 34197 24251
rect 26088 24246 34197 24248
rect 26088 24190 26093 24246
rect 26149 24190 34136 24246
rect 34192 24190 34197 24246
rect 26088 24188 34197 24190
rect 26088 24185 26154 24188
rect 34131 24185 34197 24188
rect 23256 24072 24012 24148
rect 8840 23806 8846 23870
rect 8910 23806 9052 23870
rect 8840 23800 9052 23806
rect 41616 24006 41828 24012
rect 41616 23942 41622 24006
rect 41686 23964 41828 24006
rect 41686 23942 41712 23964
rect 41616 23908 41712 23942
rect 41768 23908 41828 23964
rect 41616 23876 41828 23908
rect 41616 23870 42236 23876
rect 41616 23806 42166 23870
rect 42230 23806 42236 23870
rect 41616 23800 42236 23806
rect 34136 23598 34348 23604
rect 34136 23534 34142 23598
rect 34206 23534 34348 23598
rect 8432 23434 8644 23468
rect 8432 23378 8500 23434
rect 8556 23378 8644 23434
rect 19584 23462 24012 23468
rect 19584 23398 19726 23462
rect 19790 23398 23942 23462
rect 24006 23398 24012 23462
rect 19584 23392 24012 23398
rect 34136 23392 34348 23534
rect 39304 23528 40196 23604
rect 39304 23392 39516 23528
rect 39984 23468 40196 23528
rect 39984 23462 42916 23468
rect 39984 23398 40126 23462
rect 40190 23398 42846 23462
rect 42910 23398 42916 23462
rect 39984 23392 42916 23398
rect 8432 23332 8644 23378
rect 0 23256 8644 23332
rect 9440 23365 9506 23368
rect 9774 23365 9840 23368
rect 9440 23363 9840 23365
rect 9440 23307 9445 23363
rect 9501 23307 9779 23363
rect 9835 23307 9840 23363
rect 19709 23359 19807 23392
rect 20055 23359 20153 23392
rect 20957 23359 21055 23392
rect 21303 23359 21401 23392
rect 22205 23359 22303 23392
rect 22551 23359 22649 23392
rect 23453 23359 23551 23392
rect 23799 23359 23897 23392
rect 9440 23305 9840 23307
rect 9440 23302 9506 23305
rect 9774 23302 9840 23305
rect 40787 23096 40793 23098
rect 29158 23036 29218 23096
rect 33996 23036 40793 23096
rect 40787 23034 40793 23036
rect 40857 23034 40863 23098
rect 27897 22797 27963 22800
rect 34131 22797 34197 22800
rect 27897 22795 34197 22797
rect 27897 22739 27902 22795
rect 27958 22739 34136 22795
rect 34192 22739 34197 22795
rect 27897 22737 34197 22739
rect 27897 22734 27963 22737
rect 34131 22734 34197 22737
rect 8840 22646 9052 22652
rect 8840 22582 8982 22646
rect 9046 22582 9052 22646
rect 8840 22516 9052 22582
rect 8840 22510 12316 22516
rect 8840 22446 12246 22510
rect 12310 22446 12316 22510
rect 8840 22440 12316 22446
rect 1632 22284 1844 22380
rect 1632 22244 1730 22284
rect 1224 22238 1730 22244
rect 1224 22174 1230 22238
rect 1294 22228 1730 22238
rect 1786 22228 1844 22284
rect 1294 22174 1844 22228
rect 1224 22168 1844 22174
rect 19448 22374 19660 22380
rect 19448 22310 19590 22374
rect 19654 22310 19660 22374
rect 19448 22238 19660 22310
rect 19448 22174 19590 22238
rect 19654 22174 19660 22238
rect 19448 22168 19660 22174
rect 20264 22304 20884 22380
rect 20264 22238 20476 22304
rect 20264 22174 20270 22238
rect 20334 22174 20476 22238
rect 20264 22168 20476 22174
rect 20672 22238 20884 22304
rect 20672 22174 20814 22238
rect 20878 22174 20884 22238
rect 20672 22168 20884 22174
rect 21488 22304 22108 22380
rect 21488 22168 21700 22304
rect 21896 22238 22108 22304
rect 21896 22174 22038 22238
rect 22102 22174 22108 22238
rect 21896 22168 22108 22174
rect 22712 22304 23332 22380
rect 22712 22238 22924 22304
rect 22712 22174 22718 22238
rect 22782 22174 22924 22238
rect 22712 22168 22924 22174
rect 23120 22238 23332 22304
rect 23120 22174 23262 22238
rect 23326 22174 23332 22238
rect 23120 22168 23332 22174
rect 23936 22238 24284 22380
rect 23936 22174 24078 22238
rect 24142 22174 24284 22238
rect 23936 22168 24284 22174
rect 24344 22238 24556 22380
rect 41616 22284 41828 22380
rect 41616 22244 41712 22284
rect 24344 22174 24350 22238
rect 24414 22174 24556 22238
rect 24344 22168 24556 22174
rect 34136 22238 34348 22244
rect 34136 22174 34278 22238
rect 34342 22174 34348 22238
rect 34136 21896 34348 22174
rect 39304 22108 39516 22244
rect 39984 22228 41712 22244
rect 41768 22244 41828 22284
rect 41768 22238 42236 22244
rect 41768 22228 42166 22238
rect 39984 22174 42166 22228
rect 42230 22174 42236 22238
rect 39984 22168 42236 22174
rect 39984 22108 40196 22168
rect 39304 22032 40196 22108
rect 39304 21896 39516 22032
rect 39984 21896 40196 22032
rect 8432 21734 8644 21836
rect 9440 21807 9506 21810
rect 9694 21807 9760 21810
rect 9440 21805 9760 21807
rect 9440 21749 9445 21805
rect 9501 21749 9699 21805
rect 9755 21749 9760 21805
rect 9440 21747 9760 21749
rect 9440 21744 9506 21747
rect 9694 21744 9760 21747
rect 8432 21700 8500 21734
rect 0 21678 8500 21700
rect 8556 21678 8644 21734
rect 18904 21700 19116 21836
rect 19448 21830 20340 21836
rect 19448 21766 19590 21830
rect 19654 21766 20270 21830
rect 20334 21766 20340 21830
rect 19448 21760 20340 21766
rect 19448 21700 19796 21760
rect 18126 21694 19796 21700
rect 0 21624 8644 21678
rect 18088 21630 18094 21694
rect 18158 21630 19796 21694
rect 18126 21624 19796 21630
rect 20128 21624 20340 21760
rect 20808 21830 21020 21836
rect 20808 21766 20814 21830
rect 20878 21766 21020 21830
rect 20808 21700 21020 21766
rect 21352 21700 21564 21836
rect 22032 21830 22244 21836
rect 22032 21766 22038 21830
rect 22102 21766 22244 21830
rect 22032 21700 22244 21766
rect 22576 21830 22924 21836
rect 22576 21766 22718 21830
rect 22782 21766 22924 21830
rect 22576 21700 22924 21766
rect 20808 21624 22924 21700
rect 23256 21830 24420 21836
rect 23256 21766 23262 21830
rect 23326 21766 24078 21830
rect 24142 21766 24350 21830
rect 24414 21766 24420 21830
rect 23256 21760 24420 21766
rect 23256 21624 23468 21760
rect 23936 21700 24148 21760
rect 24480 21700 24692 21836
rect 23936 21694 26324 21700
rect 23936 21630 26254 21694
rect 26318 21630 26324 21694
rect 23936 21624 26324 21630
rect 17816 21558 19796 21564
rect 17816 21494 19726 21558
rect 19790 21494 19796 21558
rect 17816 21488 19796 21494
rect 9526 21483 9610 21487
rect 9526 21478 9643 21483
rect 9526 21422 9582 21478
rect 9638 21422 9643 21478
rect 9526 21417 9643 21422
rect 17816 21428 18028 21488
rect 9526 21413 9610 21417
rect 17816 21352 18300 21428
rect 18224 21292 18300 21352
rect 25568 21352 25780 21564
rect 26248 21422 26460 21428
rect 26248 21358 26254 21422
rect 26318 21358 26460 21422
rect 25568 21292 25644 21352
rect 8840 21286 9052 21292
rect 8840 21222 8846 21286
rect 8910 21222 9052 21286
rect 8840 21156 9052 21222
rect 3264 20884 3476 21156
rect 3944 20884 4292 21156
rect 8840 21150 10548 21156
rect 8840 21086 10478 21150
rect 10542 21086 10548 21150
rect 8840 21080 10548 21086
rect 18224 21080 18436 21292
rect 25160 21216 25644 21292
rect 26248 21292 26460 21358
rect 27200 21292 27412 21428
rect 26248 21286 27956 21292
rect 26248 21222 27886 21286
rect 27950 21222 27956 21286
rect 26248 21216 27956 21222
rect 28016 21286 28228 21428
rect 28016 21222 28022 21286
rect 28086 21222 28228 21286
rect 28016 21216 28228 21222
rect 25160 21080 25372 21216
rect 18360 21020 18436 21080
rect 25296 21020 25372 21080
rect 3264 20878 4292 20884
rect 3264 20814 3950 20878
rect 4014 20814 4292 20878
rect 3264 20808 4292 20814
rect 1632 20604 1844 20748
rect 14144 20742 14356 20884
rect 14144 20678 14150 20742
rect 14214 20678 14356 20742
rect 14144 20672 14356 20678
rect 14552 20742 14764 20884
rect 14552 20678 14694 20742
rect 14758 20678 14764 20742
rect 14552 20672 14764 20678
rect 14960 20742 15172 20884
rect 14960 20678 14966 20742
rect 15030 20678 15172 20742
rect 14960 20672 15172 20678
rect 15232 20878 18164 20884
rect 15232 20814 18094 20878
rect 18158 20814 18164 20878
rect 15232 20808 18164 20814
rect 18224 20808 18436 21020
rect 15232 20742 15580 20808
rect 18360 20748 18436 20808
rect 15232 20678 15238 20742
rect 15302 20678 15580 20742
rect 15232 20672 15580 20678
rect 1632 20548 1730 20604
rect 1786 20548 1844 20604
rect 1632 20476 1844 20548
rect 18224 20536 18436 20748
rect 25160 20808 25372 21020
rect 27918 20878 28364 20884
rect 27880 20814 27886 20878
rect 27950 20814 28022 20878
rect 28086 20814 28364 20878
rect 27918 20808 28364 20814
rect 25160 20748 25236 20808
rect 25160 20536 25372 20748
rect 28016 20742 28364 20808
rect 28016 20678 28022 20742
rect 28086 20678 28364 20742
rect 28016 20672 28364 20678
rect 28424 20742 28772 20884
rect 28424 20678 28702 20742
rect 28766 20678 28772 20742
rect 28424 20672 28772 20678
rect 28832 20742 29044 20884
rect 28832 20678 28974 20742
rect 29038 20678 29044 20742
rect 28832 20672 29044 20678
rect 29240 20742 29452 20884
rect 29240 20678 29382 20742
rect 29446 20678 29452 20742
rect 29240 20672 29452 20678
rect 39304 20612 39516 20748
rect 39984 20742 40196 20748
rect 39984 20678 40126 20742
rect 40190 20678 40196 20742
rect 39984 20612 40196 20678
rect 39304 20536 40196 20612
rect 41616 20604 41828 20748
rect 41616 20548 41712 20604
rect 41768 20548 41828 20604
rect 18224 20476 18300 20536
rect 25160 20476 25236 20536
rect 41616 20476 41828 20548
rect 1224 20470 1844 20476
rect 1224 20406 1230 20470
rect 1294 20406 1844 20470
rect 1224 20400 1844 20406
rect 14144 20470 14356 20476
rect 14144 20406 14150 20470
rect 14214 20406 14356 20470
rect 2640 20345 2706 20346
rect 2598 20281 2641 20345
rect 2705 20281 2748 20345
rect 14144 20334 14356 20406
rect 2640 20280 2706 20281
rect 14144 20270 14150 20334
rect 14214 20270 14356 20334
rect 14144 20264 14356 20270
rect 14552 20470 14764 20476
rect 14552 20406 14694 20470
rect 14758 20406 14764 20470
rect 14552 20334 14764 20406
rect 14552 20270 14694 20334
rect 14758 20270 14764 20334
rect 14552 20264 14764 20270
rect 14960 20470 15172 20476
rect 14960 20406 14966 20470
rect 15030 20406 15172 20470
rect 14960 20334 15172 20406
rect 14960 20270 14966 20334
rect 15030 20270 15172 20334
rect 14960 20264 15172 20270
rect 15232 20470 15580 20476
rect 15232 20406 15238 20470
rect 15302 20406 15580 20470
rect 15232 20334 15580 20406
rect 15232 20270 15238 20334
rect 15302 20270 15580 20334
rect 15232 20264 15580 20270
rect 18224 20264 18436 20476
rect 25160 20264 25372 20476
rect 28016 20470 28364 20476
rect 28016 20406 28022 20470
rect 28086 20406 28364 20470
rect 28016 20334 28364 20406
rect 28016 20270 28022 20334
rect 28086 20270 28364 20334
rect 28016 20264 28364 20270
rect 28424 20470 28772 20476
rect 28424 20406 28702 20470
rect 28766 20406 28772 20470
rect 28424 20334 28772 20406
rect 28424 20270 28702 20334
rect 28766 20270 28772 20334
rect 28424 20264 28772 20270
rect 28832 20470 29044 20476
rect 28832 20406 28974 20470
rect 29038 20406 29044 20470
rect 28832 20334 29044 20406
rect 28832 20270 28974 20334
rect 29038 20270 29044 20334
rect 28832 20264 29044 20270
rect 29240 20470 29452 20476
rect 29240 20406 29382 20470
rect 29446 20406 29452 20470
rect 29240 20334 29452 20406
rect 41616 20470 42236 20476
rect 41616 20406 42166 20470
rect 42230 20406 42236 20470
rect 41616 20400 42236 20406
rect 29240 20270 29246 20334
rect 29310 20270 29452 20334
rect 29240 20264 29452 20270
rect 18360 20204 18436 20264
rect 25296 20204 25372 20264
rect 14144 20062 14356 20068
rect 14144 19998 14150 20062
rect 14214 19998 14356 20062
rect 14144 19926 14356 19998
rect 14144 19862 14150 19926
rect 14214 19862 14356 19926
rect 14144 19856 14356 19862
rect 14552 20062 14764 20068
rect 14552 19998 14694 20062
rect 14758 19998 14764 20062
rect 14552 19926 14764 19998
rect 14552 19862 14558 19926
rect 14622 19862 14764 19926
rect 14552 19856 14764 19862
rect 14960 20062 15172 20068
rect 14960 19998 14966 20062
rect 15030 19998 15172 20062
rect 14960 19926 15172 19998
rect 14960 19862 15102 19926
rect 15166 19862 15172 19926
rect 14960 19856 15172 19862
rect 15232 20062 15580 20068
rect 15232 19998 15238 20062
rect 15302 19998 15580 20062
rect 15232 19926 15580 19998
rect 15232 19862 15238 19926
rect 15302 19862 15580 19926
rect 15232 19856 15580 19862
rect 18224 19992 18436 20204
rect 25160 19992 25372 20204
rect 28016 20062 28364 20068
rect 28016 19998 28022 20062
rect 28086 19998 28364 20062
rect 18224 19932 18300 19992
rect 25160 19932 25236 19992
rect 18224 19720 18436 19932
rect 18360 19660 18436 19720
rect 3264 19524 3476 19660
rect 3944 19524 4292 19660
rect 2486 19518 4292 19524
rect 2448 19454 2454 19518
rect 2518 19454 4292 19518
rect 2486 19448 4292 19454
rect 14144 19654 14356 19660
rect 14144 19590 14150 19654
rect 14214 19590 14356 19654
rect 14144 19518 14356 19590
rect 14144 19454 14150 19518
rect 14214 19454 14356 19518
rect 14144 19448 14356 19454
rect 14552 19654 14764 19660
rect 14552 19590 14558 19654
rect 14622 19590 14764 19654
rect 14552 19518 14764 19590
rect 14552 19454 14558 19518
rect 14622 19454 14764 19518
rect 14552 19448 14764 19454
rect 14960 19654 15172 19660
rect 14960 19590 15102 19654
rect 15166 19590 15172 19654
rect 14960 19518 15172 19590
rect 14960 19454 14966 19518
rect 15030 19454 15172 19518
rect 14960 19448 15172 19454
rect 15232 19654 15580 19660
rect 15232 19590 15238 19654
rect 15302 19590 15580 19654
rect 15232 19518 15580 19590
rect 15232 19454 15238 19518
rect 15302 19454 15580 19518
rect 15232 19448 15580 19454
rect 18224 19448 18436 19660
rect 25160 19720 25372 19932
rect 28016 19926 28364 19998
rect 28016 19862 28294 19926
rect 28358 19862 28364 19926
rect 28016 19856 28364 19862
rect 28424 20062 28772 20068
rect 28424 19998 28702 20062
rect 28766 19998 28772 20062
rect 28424 19926 28772 19998
rect 28424 19862 28430 19926
rect 28494 19862 28772 19926
rect 28424 19856 28772 19862
rect 28832 20062 29044 20068
rect 28832 19998 28974 20062
rect 29038 19998 29044 20062
rect 28832 19926 29044 19998
rect 28832 19862 28838 19926
rect 28902 19862 29044 19926
rect 28832 19856 29044 19862
rect 29240 20062 29452 20068
rect 29240 19998 29246 20062
rect 29310 19998 29452 20062
rect 29240 19926 29452 19998
rect 29240 19862 29246 19926
rect 29310 19862 29452 19926
rect 29240 19856 29452 19862
rect 25160 19660 25236 19720
rect 25160 19448 25372 19660
rect 28016 19654 28364 19660
rect 28016 19590 28294 19654
rect 28358 19590 28364 19654
rect 28016 19518 28364 19590
rect 28016 19454 28158 19518
rect 28222 19454 28364 19518
rect 28016 19448 28364 19454
rect 28424 19654 28772 19660
rect 28424 19590 28430 19654
rect 28494 19590 28772 19654
rect 28424 19518 28772 19590
rect 28424 19454 28430 19518
rect 28494 19454 28772 19518
rect 28424 19448 28772 19454
rect 28832 19654 29044 19660
rect 28832 19590 28838 19654
rect 28902 19590 29044 19654
rect 28832 19518 29044 19590
rect 28832 19454 28838 19518
rect 28902 19454 29044 19518
rect 28832 19448 29044 19454
rect 29240 19654 29452 19660
rect 29240 19590 29246 19654
rect 29310 19590 29452 19654
rect 29240 19518 29452 19590
rect 29240 19454 29246 19518
rect 29310 19454 29452 19518
rect 29240 19448 29452 19454
rect 18224 19388 18300 19448
rect 25160 19388 25236 19448
rect 14144 19246 14356 19252
rect 14144 19182 14150 19246
rect 14214 19182 14356 19246
rect 14144 19040 14356 19182
rect 14552 19246 14764 19252
rect 14552 19182 14558 19246
rect 14622 19182 14764 19246
rect 14552 19040 14764 19182
rect 14960 19246 15172 19252
rect 14960 19182 14966 19246
rect 15030 19182 15172 19246
rect 14960 19110 15172 19182
rect 14960 19046 14966 19110
rect 15030 19046 15172 19110
rect 14960 19040 15172 19046
rect 15232 19246 15580 19252
rect 15232 19182 15238 19246
rect 15302 19182 15580 19246
rect 15232 19110 15580 19182
rect 18224 19176 18436 19388
rect 25160 19176 25372 19388
rect 39304 19312 40196 19388
rect 18360 19116 18436 19176
rect 25296 19116 25372 19176
rect 15232 19046 15238 19110
rect 15302 19046 15580 19110
rect 15232 19040 15580 19046
rect 14144 18980 14220 19040
rect 14552 18980 14628 19040
rect 1224 18974 2524 18980
rect 1224 18910 1230 18974
rect 1294 18924 2454 18974
rect 1294 18910 1730 18924
rect 1224 18904 1730 18910
rect 1632 18868 1730 18904
rect 1786 18910 2454 18924
rect 2518 18910 2524 18974
rect 1786 18904 2524 18910
rect 1786 18868 1844 18904
rect 1632 18768 1844 18868
rect 14144 18632 14356 18980
rect 14552 18632 14764 18980
rect 18224 18904 18436 19116
rect 25160 18974 25372 19116
rect 28016 19246 28364 19252
rect 28016 19182 28158 19246
rect 28222 19182 28364 19246
rect 28016 19110 28364 19182
rect 28016 19046 28022 19110
rect 28086 19046 28364 19110
rect 28016 19040 28364 19046
rect 28424 19246 28772 19252
rect 28424 19182 28430 19246
rect 28494 19182 28772 19246
rect 28424 19110 28772 19182
rect 28424 19046 28430 19110
rect 28494 19046 28772 19110
rect 28424 19040 28772 19046
rect 28832 19246 29044 19252
rect 28832 19182 28838 19246
rect 28902 19182 29044 19246
rect 28832 19040 29044 19182
rect 28968 18980 29044 19040
rect 25160 18910 25166 18974
rect 25230 18910 25372 18974
rect 25160 18904 25372 18910
rect 18224 18844 18300 18904
rect 25296 18844 25372 18904
rect 14960 18838 15172 18844
rect 14960 18774 14966 18838
rect 15030 18774 15172 18838
rect 14960 18702 15172 18774
rect 14960 18638 15102 18702
rect 15166 18638 15172 18702
rect 14960 18632 15172 18638
rect 15232 18838 15580 18844
rect 15232 18774 15238 18838
rect 15302 18774 15580 18838
rect 15232 18702 15580 18774
rect 15232 18638 15374 18702
rect 15438 18638 15580 18702
rect 15232 18632 15580 18638
rect 14144 18572 14220 18632
rect 14552 18572 14628 18632
rect 11696 18300 12044 18572
rect 12240 18566 12996 18572
rect 12240 18502 12246 18566
rect 12310 18502 12996 18566
rect 12240 18496 12996 18502
rect 3264 18294 4292 18300
rect 3264 18230 3950 18294
rect 4014 18230 4292 18294
rect 3264 18224 4292 18230
rect 11696 18294 12180 18300
rect 11696 18230 11838 18294
rect 11902 18230 12180 18294
rect 11696 18224 12180 18230
rect 12240 18294 12452 18496
rect 12920 18436 12996 18496
rect 12240 18230 12246 18294
rect 12310 18230 12382 18294
rect 12446 18230 12452 18294
rect 12240 18224 12452 18230
rect 12512 18294 12860 18436
rect 12512 18230 12518 18294
rect 12582 18230 12860 18294
rect 12512 18224 12860 18230
rect 12920 18224 13132 18436
rect 14144 18224 14356 18572
rect 14552 18224 14764 18572
rect 15096 18566 15852 18572
rect 15096 18502 15782 18566
rect 15846 18502 15852 18566
rect 15096 18496 15852 18502
rect 15096 18436 15172 18496
rect 14960 18430 15172 18436
rect 14960 18366 15102 18430
rect 15166 18366 15172 18430
rect 14960 18224 15172 18366
rect 15232 18430 15580 18436
rect 15232 18366 15374 18430
rect 15438 18366 15580 18430
rect 15232 18300 15580 18366
rect 18224 18430 18436 18844
rect 18224 18366 18230 18430
rect 18294 18366 18436 18430
rect 18224 18360 18436 18366
rect 18360 18300 18436 18360
rect 15232 18294 16260 18300
rect 15232 18230 16190 18294
rect 16254 18230 16260 18294
rect 15232 18224 16260 18230
rect 17000 18224 18164 18300
rect 3264 18164 3476 18224
rect 544 18158 3884 18164
rect 544 18094 550 18158
rect 614 18094 3814 18158
rect 3878 18094 3884 18158
rect 544 18088 3884 18094
rect 3944 18088 4292 18224
rect 12104 18164 12180 18224
rect 12512 18164 12588 18224
rect 12104 18088 12588 18164
rect 14144 18164 14220 18224
rect 14552 18164 14628 18224
rect 14960 18164 15036 18224
rect 15232 18164 15308 18224
rect 17000 18164 17076 18224
rect 18088 18164 18164 18224
rect 18224 18164 18436 18300
rect 14144 18022 14356 18164
rect 14144 17958 14150 18022
rect 14214 17958 14356 18022
rect 14144 17952 14356 17958
rect 14552 18022 14764 18164
rect 14552 17958 14694 18022
rect 14758 17958 14764 18022
rect 14552 17952 14764 17958
rect 10744 17816 11772 17892
rect 10744 17756 10820 17816
rect 11696 17756 11772 17816
rect 12376 17816 12996 17892
rect 12376 17756 12452 17816
rect 12920 17756 12996 17816
rect 14960 17816 15172 18164
rect 15232 17816 15580 18164
rect 16048 18088 17076 18164
rect 16048 18028 16124 18088
rect 15776 18022 16124 18028
rect 15776 17958 15782 18022
rect 15846 17958 16124 18022
rect 15776 17952 16124 17958
rect 16184 18022 16396 18028
rect 16184 17958 16190 18022
rect 16254 17958 16396 18022
rect 15776 17816 15988 17952
rect 16184 17892 16396 17958
rect 16184 17816 16532 17892
rect 16592 17816 16804 18088
rect 17136 17816 17484 18164
rect 18088 18158 18436 18164
rect 18088 18094 18230 18158
rect 18294 18094 18436 18158
rect 18088 18088 18436 18094
rect 14960 17756 15036 17816
rect 15232 17756 15308 17816
rect 16456 17756 16532 17816
rect 17136 17756 17212 17816
rect 10472 17750 10820 17756
rect 10472 17686 10478 17750
rect 10542 17686 10820 17750
rect 10472 17680 10820 17686
rect 10472 17408 10684 17680
rect 10880 17484 11092 17756
rect 11696 17750 12044 17756
rect 11696 17686 11838 17750
rect 11902 17686 12044 17750
rect 11696 17544 12044 17686
rect 12240 17750 12452 17756
rect 12240 17686 12382 17750
rect 12446 17686 12452 17750
rect 12240 17544 12452 17686
rect 12512 17750 12860 17756
rect 12512 17686 12518 17750
rect 12582 17686 12860 17750
rect 10880 17478 12316 17484
rect 10880 17414 12246 17478
rect 12310 17414 12316 17478
rect 10880 17408 12316 17414
rect 12512 17478 12860 17686
rect 12512 17414 12654 17478
rect 12718 17414 12860 17478
rect 12512 17408 12860 17414
rect 12920 17478 13132 17756
rect 14144 17750 14356 17756
rect 14144 17686 14150 17750
rect 14214 17686 14356 17750
rect 14144 17614 14356 17686
rect 14144 17550 14150 17614
rect 14214 17550 14356 17614
rect 14144 17544 14356 17550
rect 14552 17750 14764 17756
rect 14552 17686 14694 17750
rect 14758 17686 14764 17750
rect 14552 17614 14764 17686
rect 14552 17550 14694 17614
rect 14758 17550 14764 17614
rect 14552 17544 14764 17550
rect 14960 17484 15172 17756
rect 12920 17414 13062 17478
rect 13126 17414 13132 17478
rect 12920 17408 13132 17414
rect 14416 17408 15172 17484
rect 14416 17348 14492 17408
rect 15096 17348 15172 17408
rect 1632 17244 1844 17348
rect 1632 17212 1730 17244
rect 1224 17206 1730 17212
rect 1224 17142 1230 17206
rect 1294 17188 1730 17206
rect 1786 17212 1844 17244
rect 14144 17342 14492 17348
rect 14144 17278 14150 17342
rect 14214 17278 14492 17342
rect 14144 17272 14492 17278
rect 14552 17342 14764 17348
rect 14552 17278 14694 17342
rect 14758 17278 14764 17342
rect 1786 17206 3340 17212
rect 1786 17188 3270 17206
rect 1294 17142 3270 17188
rect 3334 17142 3340 17206
rect 1224 17136 3340 17142
rect 14144 17206 14356 17272
rect 14144 17142 14286 17206
rect 14350 17142 14356 17206
rect 14144 17136 14356 17142
rect 14552 17206 14764 17278
rect 14552 17142 14694 17206
rect 14758 17142 14764 17206
rect 14552 17136 14764 17142
rect 14960 17206 15172 17348
rect 14960 17142 15102 17206
rect 15166 17142 15172 17206
rect 14960 17136 15172 17142
rect 15232 17408 15580 17756
rect 16456 17680 17212 17756
rect 18224 17750 18436 18088
rect 18224 17686 18366 17750
rect 18430 17686 18436 17750
rect 18224 17680 18436 17686
rect 25160 18702 25372 18844
rect 25160 18638 25166 18702
rect 25230 18638 25372 18702
rect 25160 18360 25372 18638
rect 28016 18838 28364 18844
rect 28016 18774 28022 18838
rect 28086 18774 28364 18838
rect 28016 18702 28364 18774
rect 28016 18638 28158 18702
rect 28222 18638 28364 18702
rect 28016 18632 28364 18638
rect 28424 18838 28772 18844
rect 28424 18774 28430 18838
rect 28494 18774 28772 18838
rect 28424 18702 28772 18774
rect 28424 18638 28702 18702
rect 28766 18638 28772 18702
rect 28424 18632 28772 18638
rect 28832 18632 29044 18980
rect 28968 18572 29044 18632
rect 27918 18566 28500 18572
rect 27880 18502 27886 18566
rect 27950 18502 28500 18566
rect 27918 18496 28500 18502
rect 28424 18436 28500 18496
rect 28016 18430 28364 18436
rect 28016 18366 28158 18430
rect 28222 18366 28364 18430
rect 25160 18300 25236 18360
rect 25160 17756 25372 18300
rect 27336 18294 27684 18300
rect 27336 18230 27614 18294
rect 27678 18230 27684 18294
rect 27336 18224 27684 18230
rect 28016 18224 28364 18366
rect 28424 18430 28772 18436
rect 28424 18366 28702 18430
rect 28766 18366 28772 18430
rect 28424 18224 28772 18366
rect 28832 18224 29044 18572
rect 29240 19246 29452 19252
rect 29240 19182 29246 19246
rect 29310 19182 29452 19246
rect 29240 19040 29452 19182
rect 39304 19176 39516 19312
rect 39984 19252 40196 19312
rect 39984 19246 41692 19252
rect 39984 19182 41622 19246
rect 41686 19182 41692 19246
rect 39984 19176 41692 19182
rect 29240 18980 29316 19040
rect 29240 18632 29452 18980
rect 41616 18974 42236 18980
rect 41616 18910 41622 18974
rect 41686 18924 42166 18974
rect 41686 18910 41712 18924
rect 41616 18868 41712 18910
rect 41768 18910 42166 18924
rect 42230 18910 42236 18974
rect 41768 18904 42236 18910
rect 41768 18868 41828 18904
rect 41616 18768 41828 18868
rect 29240 18572 29316 18632
rect 29240 18224 29452 18572
rect 30736 18496 31492 18572
rect 30736 18436 30812 18496
rect 30464 18360 30812 18436
rect 30464 18294 30676 18360
rect 30464 18230 30470 18294
rect 30534 18230 30676 18294
rect 30464 18224 30676 18230
rect 30872 18224 31084 18436
rect 31144 18294 31492 18496
rect 31144 18230 31150 18294
rect 31214 18230 31492 18294
rect 31144 18224 31492 18230
rect 31552 18294 31900 18572
rect 31552 18230 31694 18294
rect 31758 18230 31900 18294
rect 31552 18224 31900 18230
rect 27336 18164 27412 18224
rect 28152 18164 28228 18224
rect 28560 18164 28636 18224
rect 28832 18164 28908 18224
rect 29240 18164 29316 18224
rect 31008 18164 31084 18224
rect 31552 18164 31628 18224
rect 26248 17892 26460 18164
rect 26792 18088 27412 18164
rect 27472 18088 28364 18164
rect 26792 18028 27004 18088
rect 27472 18028 27548 18088
rect 26558 18022 27004 18028
rect 26520 17958 26526 18022
rect 26590 17958 27004 18022
rect 26558 17952 27004 17958
rect 26248 17816 26732 17892
rect 26792 17816 27004 17952
rect 27200 17952 27548 18028
rect 27608 18022 27956 18028
rect 27608 17958 27614 18022
rect 27678 17958 27886 18022
rect 27950 17958 27956 18022
rect 27608 17952 27956 17958
rect 27200 17816 27412 17952
rect 27608 17816 27820 17952
rect 28016 17816 28364 18088
rect 28424 17892 28772 18164
rect 28832 18022 29044 18164
rect 28832 17958 28974 18022
rect 29038 17958 29044 18022
rect 28832 17952 29044 17958
rect 29240 18022 29452 18164
rect 31008 18088 31628 18164
rect 29240 17958 29246 18022
rect 29310 17958 29452 18022
rect 29240 17952 29452 17958
rect 28424 17816 29316 17892
rect 26656 17756 26732 17816
rect 27200 17756 27276 17816
rect 28288 17756 28364 17816
rect 28560 17756 28636 17816
rect 29240 17756 29316 17816
rect 31008 17816 31628 17892
rect 31008 17756 31084 17816
rect 31552 17756 31628 17816
rect 32368 17816 32988 17892
rect 32368 17756 32444 17816
rect 32912 17756 32988 17816
rect 39304 17886 42916 17892
rect 39304 17822 42846 17886
rect 42910 17822 42916 17886
rect 39304 17816 42916 17822
rect 25160 17750 26596 17756
rect 25160 17686 25302 17750
rect 25366 17686 26526 17750
rect 26590 17686 26596 17750
rect 25160 17680 26596 17686
rect 26656 17680 27276 17756
rect 18224 17478 18436 17484
rect 18224 17414 18366 17478
rect 18430 17414 18436 17478
rect 15232 17348 15308 17408
rect 15232 17206 15580 17348
rect 15232 17142 15238 17206
rect 15302 17142 15580 17206
rect 15232 17136 15580 17142
rect 18224 17342 18436 17414
rect 18224 17278 18366 17342
rect 18430 17278 18436 17342
rect 18224 17136 18436 17278
rect 25160 17478 25372 17484
rect 25160 17414 25302 17478
rect 25366 17414 25372 17478
rect 25160 17342 25372 17414
rect 28016 17408 28364 17756
rect 28424 17408 28772 17756
rect 28832 17750 29044 17756
rect 28832 17686 28974 17750
rect 29038 17686 29044 17750
rect 28832 17614 29044 17686
rect 28832 17550 28974 17614
rect 29038 17550 29044 17614
rect 28832 17544 29044 17550
rect 29240 17750 29452 17756
rect 29240 17686 29246 17750
rect 29310 17686 29452 17750
rect 29240 17614 29452 17686
rect 29240 17550 29246 17614
rect 29310 17550 29452 17614
rect 29240 17544 29452 17550
rect 30464 17750 30676 17756
rect 30464 17686 30470 17750
rect 30534 17686 30676 17750
rect 30464 17478 30676 17686
rect 30464 17414 30470 17478
rect 30534 17414 30676 17478
rect 30464 17408 30676 17414
rect 30872 17478 31084 17756
rect 31144 17750 31492 17756
rect 31144 17686 31150 17750
rect 31214 17686 31492 17750
rect 31144 17544 31492 17686
rect 31552 17750 32444 17756
rect 31552 17686 31694 17750
rect 31758 17686 32444 17750
rect 31552 17680 32444 17686
rect 31552 17544 31900 17680
rect 30872 17414 30878 17478
rect 30942 17414 31084 17478
rect 30872 17408 31084 17414
rect 31416 17484 31492 17544
rect 32504 17484 32716 17756
rect 31416 17408 32716 17484
rect 32912 17408 33124 17756
rect 39304 17680 39516 17816
rect 39984 17756 40196 17816
rect 39886 17750 40196 17756
rect 39848 17686 39854 17750
rect 39918 17686 40196 17750
rect 39886 17680 40196 17686
rect 28152 17348 28228 17408
rect 28696 17348 28772 17408
rect 25160 17278 25302 17342
rect 25366 17278 25372 17342
rect 25160 17136 25372 17278
rect 28016 17206 28364 17348
rect 28016 17142 28158 17206
rect 28222 17142 28364 17206
rect 28016 17136 28364 17142
rect 28424 17206 28772 17348
rect 28424 17142 28702 17206
rect 28766 17142 28772 17206
rect 28424 17136 28772 17142
rect 28832 17342 29044 17348
rect 28832 17278 28974 17342
rect 29038 17278 29044 17342
rect 28832 17206 29044 17278
rect 28832 17142 28974 17206
rect 29038 17142 29044 17206
rect 28832 17136 29044 17142
rect 29240 17342 29452 17348
rect 29240 17278 29246 17342
rect 29310 17278 29452 17342
rect 29240 17206 29452 17278
rect 29240 17142 29246 17206
rect 29310 17142 29452 17206
rect 29240 17136 29452 17142
rect 41616 17244 41828 17348
rect 41616 17206 41712 17244
rect 41616 17142 41622 17206
rect 41686 17188 41712 17206
rect 41768 17212 41828 17244
rect 41768 17206 42236 17212
rect 41768 17188 42166 17206
rect 41686 17142 42166 17188
rect 42230 17142 42236 17206
rect 41616 17136 42236 17142
rect 18360 17076 18436 17136
rect 25296 17076 25372 17136
rect 18224 17070 18436 17076
rect 18224 17006 18366 17070
rect 18430 17006 18436 17070
rect 14144 16934 14356 16940
rect 14144 16870 14286 16934
rect 14350 16870 14356 16934
rect 3264 16798 4292 16804
rect 3264 16734 3270 16798
rect 3334 16734 4292 16798
rect 3264 16728 4292 16734
rect 14144 16798 14356 16870
rect 14144 16734 14150 16798
rect 14214 16734 14356 16798
rect 14144 16728 14356 16734
rect 14552 16934 14764 16940
rect 14552 16870 14694 16934
rect 14758 16870 14764 16934
rect 14552 16798 14764 16870
rect 14552 16734 14558 16798
rect 14622 16734 14764 16798
rect 14552 16728 14764 16734
rect 14960 16934 15172 16940
rect 14960 16870 15102 16934
rect 15166 16870 15172 16934
rect 14960 16798 15172 16870
rect 14960 16734 15102 16798
rect 15166 16734 15172 16798
rect 14960 16728 15172 16734
rect 15232 16934 15580 16940
rect 15232 16870 15238 16934
rect 15302 16870 15580 16934
rect 15232 16798 15580 16870
rect 18224 16864 18436 17006
rect 25160 17070 25372 17076
rect 25160 17006 25302 17070
rect 25366 17006 25372 17070
rect 25160 16864 25372 17006
rect 18360 16804 18436 16864
rect 25296 16804 25372 16864
rect 15232 16734 15510 16798
rect 15574 16734 15580 16798
rect 15232 16728 15580 16734
rect 3264 16592 3476 16728
rect 3944 16592 4292 16728
rect 18224 16592 18436 16804
rect 18360 16532 18436 16592
rect 14144 16526 14356 16532
rect 14144 16462 14150 16526
rect 14214 16462 14356 16526
rect 14144 16390 14356 16462
rect 14144 16326 14286 16390
rect 14350 16326 14356 16390
rect 14144 16320 14356 16326
rect 14552 16526 14764 16532
rect 14552 16462 14558 16526
rect 14622 16462 14764 16526
rect 14552 16390 14764 16462
rect 14552 16326 14694 16390
rect 14758 16326 14764 16390
rect 14552 16320 14764 16326
rect 14960 16526 15172 16532
rect 14960 16462 15102 16526
rect 15166 16462 15172 16526
rect 14960 16390 15172 16462
rect 14960 16326 15102 16390
rect 15166 16326 15172 16390
rect 14960 16320 15172 16326
rect 15232 16526 15580 16532
rect 15232 16462 15510 16526
rect 15574 16462 15580 16526
rect 15232 16390 15580 16462
rect 15232 16326 15510 16390
rect 15574 16326 15580 16390
rect 15232 16320 15580 16326
rect 18224 16320 18436 16532
rect 25160 16592 25372 16804
rect 28016 16934 28364 16940
rect 28016 16870 28158 16934
rect 28222 16870 28364 16934
rect 28016 16798 28364 16870
rect 28016 16734 28158 16798
rect 28222 16734 28364 16798
rect 28016 16728 28364 16734
rect 28424 16934 28772 16940
rect 28424 16870 28702 16934
rect 28766 16870 28772 16934
rect 28424 16798 28772 16870
rect 28424 16734 28566 16798
rect 28630 16734 28772 16798
rect 28424 16728 28772 16734
rect 28832 16934 29044 16940
rect 28832 16870 28974 16934
rect 29038 16870 29044 16934
rect 28832 16798 29044 16870
rect 28832 16734 28974 16798
rect 29038 16734 29044 16798
rect 28832 16728 29044 16734
rect 29240 16934 29452 16940
rect 29240 16870 29246 16934
rect 29310 16870 29452 16934
rect 29240 16798 29452 16870
rect 29240 16734 29246 16798
rect 29310 16734 29452 16798
rect 29240 16728 29452 16734
rect 25160 16532 25236 16592
rect 25160 16320 25372 16532
rect 28016 16526 28364 16532
rect 28016 16462 28158 16526
rect 28222 16462 28364 16526
rect 28016 16390 28364 16462
rect 28016 16326 28294 16390
rect 28358 16326 28364 16390
rect 28016 16320 28364 16326
rect 28424 16526 28772 16532
rect 28424 16462 28566 16526
rect 28630 16462 28772 16526
rect 28424 16390 28772 16462
rect 28424 16326 28566 16390
rect 28630 16326 28772 16390
rect 28424 16320 28772 16326
rect 28832 16526 29044 16532
rect 28832 16462 28974 16526
rect 29038 16462 29044 16526
rect 28832 16390 29044 16462
rect 28832 16326 28974 16390
rect 29038 16326 29044 16390
rect 28832 16320 29044 16326
rect 29240 16526 29452 16532
rect 29240 16462 29246 16526
rect 29310 16462 29452 16526
rect 29240 16390 29452 16462
rect 29240 16326 29246 16390
rect 29310 16326 29452 16390
rect 29240 16320 29452 16326
rect 39304 16526 41692 16532
rect 39304 16462 41622 16526
rect 41686 16462 41692 16526
rect 39304 16456 41692 16462
rect 39304 16320 39516 16456
rect 39984 16320 40196 16456
rect 18224 16260 18300 16320
rect 25296 16260 25372 16320
rect 12376 16184 12996 16260
rect 12376 16124 12452 16184
rect 12920 16124 12996 16184
rect 11696 15988 12044 16124
rect 11696 15982 12180 15988
rect 11696 15918 11974 15982
rect 12038 15918 12180 15982
rect 11696 15912 12180 15918
rect 12240 15982 12452 16124
rect 12240 15918 12246 15982
rect 12310 15918 12452 15982
rect 12240 15912 12452 15918
rect 12512 16118 12860 16124
rect 12512 16054 12654 16118
rect 12718 16054 12860 16118
rect 12512 15982 12860 16054
rect 12512 15918 12790 15982
rect 12854 15918 12860 15982
rect 12512 15912 12860 15918
rect 12920 16118 13132 16124
rect 12920 16054 13062 16118
rect 13126 16054 13132 16118
rect 12920 15988 13132 16054
rect 14144 16118 14356 16124
rect 14144 16054 14286 16118
rect 14350 16054 14356 16118
rect 12920 15912 14084 15988
rect 14144 15982 14356 16054
rect 14144 15918 14286 15982
rect 14350 15918 14356 15982
rect 14144 15912 14356 15918
rect 14552 16118 14764 16124
rect 14552 16054 14694 16118
rect 14758 16054 14764 16118
rect 14552 15988 14764 16054
rect 14960 16118 15172 16124
rect 14960 16054 15102 16118
rect 15166 16054 15172 16118
rect 14552 15982 14900 15988
rect 14552 15918 14694 15982
rect 14758 15918 14900 15982
rect 14552 15912 14900 15918
rect 14960 15982 15172 16054
rect 14960 15918 14966 15982
rect 15030 15918 15172 15982
rect 14960 15912 15172 15918
rect 15232 16118 15580 16124
rect 15232 16054 15510 16118
rect 15574 16054 15580 16118
rect 15232 15982 15580 16054
rect 18224 16048 18436 16260
rect 25160 16048 25372 16260
rect 30328 16184 30948 16260
rect 30328 16124 30404 16184
rect 30872 16124 30948 16184
rect 31008 16184 31628 16260
rect 31008 16124 31084 16184
rect 31552 16124 31628 16184
rect 18360 15988 18436 16048
rect 25296 15988 25372 16048
rect 15232 15918 15510 15982
rect 15574 15918 15580 15982
rect 15232 15912 15580 15918
rect 12104 15852 12180 15912
rect 12512 15852 12588 15912
rect 12104 15776 12588 15852
rect 14008 15852 14084 15912
rect 14552 15852 14628 15912
rect 14008 15776 14628 15852
rect 14824 15852 14900 15912
rect 14824 15776 15308 15852
rect 15232 15716 15308 15776
rect 18224 15776 18436 15988
rect 25160 15776 25372 15988
rect 28016 16118 28364 16124
rect 28016 16054 28294 16118
rect 28358 16054 28364 16118
rect 28016 15982 28364 16054
rect 28016 15918 28158 15982
rect 28222 15918 28364 15982
rect 28016 15912 28364 15918
rect 28424 16118 28772 16124
rect 28424 16054 28566 16118
rect 28630 16054 28772 16118
rect 28424 15982 28772 16054
rect 28424 15918 28566 15982
rect 28630 15918 28772 15982
rect 28424 15912 28772 15918
rect 28832 16118 29044 16124
rect 28832 16054 28974 16118
rect 29038 16054 29044 16118
rect 28832 15988 29044 16054
rect 29240 16118 30404 16124
rect 29240 16054 29246 16118
rect 29310 16054 30404 16118
rect 29240 16048 30404 16054
rect 30464 16118 30676 16124
rect 30464 16054 30470 16118
rect 30534 16054 30676 16118
rect 28832 15982 29180 15988
rect 28832 15918 28974 15982
rect 29038 15918 29180 15982
rect 28832 15912 29180 15918
rect 29240 15982 29452 16048
rect 29240 15918 29382 15982
rect 29446 15918 29452 15982
rect 29240 15912 29452 15918
rect 30464 15988 30676 16054
rect 30872 16118 31084 16124
rect 30872 16054 30878 16118
rect 30942 16054 31084 16118
rect 30464 15912 30812 15988
rect 30872 15982 31084 16054
rect 30872 15918 31014 15982
rect 31078 15918 31084 15982
rect 30872 15912 31084 15918
rect 31144 15982 31492 16124
rect 31144 15918 31286 15982
rect 31350 15918 31492 15982
rect 31144 15912 31492 15918
rect 31552 15912 31900 16124
rect 29104 15852 29180 15912
rect 30464 15852 30540 15912
rect 29104 15776 30540 15852
rect 30736 15852 30812 15912
rect 31144 15852 31220 15912
rect 30736 15776 31220 15852
rect 18224 15716 18300 15776
rect 25296 15716 25372 15776
rect 1632 15580 1844 15716
rect 12822 15710 14356 15716
rect 12784 15646 12790 15710
rect 12854 15646 14286 15710
rect 14350 15646 14356 15710
rect 12822 15640 14356 15646
rect 1224 15574 1844 15580
rect 1224 15510 1230 15574
rect 1294 15564 1844 15574
rect 1294 15510 1730 15564
rect 1224 15508 1730 15510
rect 1786 15508 1844 15564
rect 1224 15504 1844 15508
rect 14144 15574 14356 15640
rect 14144 15510 14150 15574
rect 14214 15510 14356 15574
rect 14144 15504 14356 15510
rect 14552 15710 14764 15716
rect 14552 15646 14694 15710
rect 14758 15646 14764 15710
rect 14552 15574 14764 15646
rect 14552 15510 14694 15574
rect 14758 15510 14764 15574
rect 14552 15504 14764 15510
rect 14960 15710 15172 15716
rect 14960 15646 14966 15710
rect 15030 15646 15172 15710
rect 14960 15574 15172 15646
rect 14960 15510 14966 15574
rect 15030 15510 15172 15574
rect 14960 15504 15172 15510
rect 15232 15710 15580 15716
rect 15232 15646 15510 15710
rect 15574 15646 15580 15710
rect 15232 15574 15580 15646
rect 15232 15510 15238 15574
rect 15302 15510 15580 15574
rect 15232 15504 15580 15510
rect 18224 15504 18436 15716
rect 25160 15504 25372 15716
rect 28016 15710 28364 15716
rect 28016 15646 28158 15710
rect 28222 15646 28364 15710
rect 28016 15574 28364 15646
rect 28016 15510 28022 15574
rect 28086 15510 28364 15574
rect 28016 15504 28364 15510
rect 28424 15710 28772 15716
rect 28424 15646 28566 15710
rect 28630 15646 28772 15710
rect 28424 15574 28772 15646
rect 28424 15510 28566 15574
rect 28630 15510 28772 15574
rect 28424 15504 28772 15510
rect 28832 15710 29044 15716
rect 28832 15646 28974 15710
rect 29038 15646 29044 15710
rect 28832 15574 29044 15646
rect 28832 15510 28974 15574
rect 29038 15510 29044 15574
rect 28832 15504 29044 15510
rect 29240 15710 29452 15716
rect 29240 15646 29382 15710
rect 29446 15646 29452 15710
rect 29240 15574 29452 15646
rect 29240 15510 29246 15574
rect 29310 15510 29452 15574
rect 29240 15504 29452 15510
rect 41616 15564 41828 15716
rect 41616 15508 41712 15564
rect 41768 15508 41828 15564
rect 1632 15368 1844 15504
rect 18224 15444 18300 15504
rect 25160 15444 25236 15504
rect 41616 15444 41828 15508
rect 3264 15308 3476 15444
rect 3846 15438 4292 15444
rect 3808 15374 3814 15438
rect 3878 15374 4292 15438
rect 3846 15368 4292 15374
rect 3944 15308 4292 15368
rect 11560 15368 12316 15444
rect 11560 15308 11636 15368
rect 12240 15308 12316 15368
rect 3264 15302 4292 15308
rect 3264 15238 3406 15302
rect 3470 15238 4292 15302
rect 3264 15232 4292 15238
rect 10472 15172 10684 15308
rect 10880 15232 11636 15308
rect 11696 15302 12044 15308
rect 11696 15238 11974 15302
rect 12038 15238 12044 15302
rect 10472 15166 10820 15172
rect 10472 15102 10478 15166
rect 10542 15102 10820 15166
rect 10472 15096 10820 15102
rect 10880 15166 11092 15232
rect 10880 15102 10886 15166
rect 10950 15102 11092 15166
rect 10880 15096 11092 15102
rect 11696 15172 12044 15238
rect 12240 15302 12452 15308
rect 12240 15238 12246 15302
rect 12310 15238 12452 15302
rect 11696 15166 12180 15172
rect 11696 15102 12110 15166
rect 12174 15102 12180 15166
rect 11696 15096 12180 15102
rect 12240 15096 12452 15238
rect 12512 15166 12860 15308
rect 12512 15102 12518 15166
rect 12582 15102 12860 15166
rect 12512 15096 12860 15102
rect 12920 15096 13132 15308
rect 14144 15302 14356 15308
rect 14144 15238 14150 15302
rect 14214 15238 14356 15302
rect 14144 15096 14356 15238
rect 14552 15302 14764 15308
rect 14552 15238 14694 15302
rect 14758 15238 14764 15302
rect 14552 15096 14764 15238
rect 14960 15302 15172 15308
rect 14960 15238 14966 15302
rect 15030 15238 15172 15302
rect 14960 15096 15172 15238
rect 15232 15302 15580 15308
rect 15232 15238 15238 15302
rect 15302 15238 15580 15302
rect 15232 15166 15580 15238
rect 18224 15232 18436 15444
rect 18360 15172 18436 15232
rect 15232 15102 15374 15166
rect 15438 15102 15580 15166
rect 15232 15096 15580 15102
rect 10744 15036 10820 15096
rect 11696 15036 11772 15096
rect 10744 14960 11772 15036
rect 12376 15036 12452 15096
rect 12920 15036 12996 15096
rect 12376 14960 12996 15036
rect 18224 15030 18436 15172
rect 18224 14966 18230 15030
rect 18294 14966 18436 15030
rect 18224 14960 18436 14966
rect 18360 14900 18436 14960
rect 12142 14894 12588 14900
rect 12104 14830 12110 14894
rect 12174 14830 12518 14894
rect 12582 14830 12588 14894
rect 12142 14824 12588 14830
rect 18224 14764 18436 14900
rect 25160 15232 25372 15444
rect 31008 15368 31628 15444
rect 31008 15308 31084 15368
rect 31552 15308 31628 15368
rect 32368 15368 32988 15444
rect 41616 15438 42236 15444
rect 41616 15374 42166 15438
rect 42230 15374 42236 15438
rect 41616 15368 42236 15374
rect 32368 15308 32444 15368
rect 32912 15308 32988 15368
rect 28016 15302 28364 15308
rect 28016 15238 28022 15302
rect 28086 15238 28364 15302
rect 25160 15172 25236 15232
rect 25160 14960 25372 15172
rect 28016 15096 28364 15238
rect 28424 15302 28772 15308
rect 28424 15238 28566 15302
rect 28630 15238 28772 15302
rect 28424 15096 28772 15238
rect 28832 15302 29044 15308
rect 28832 15238 28974 15302
rect 29038 15238 29044 15302
rect 28832 15096 29044 15238
rect 29240 15302 29452 15308
rect 29240 15238 29246 15302
rect 29310 15238 29452 15302
rect 29240 15096 29452 15238
rect 30464 15172 30676 15308
rect 30872 15302 31084 15308
rect 30872 15238 31014 15302
rect 31078 15238 31084 15302
rect 30464 15096 30812 15172
rect 30872 15096 31084 15238
rect 31144 15302 31492 15308
rect 31144 15238 31286 15302
rect 31350 15238 31492 15302
rect 31144 15096 31492 15238
rect 31552 15232 32444 15308
rect 31552 15096 31900 15232
rect 32504 15172 32716 15308
rect 32912 15172 33124 15308
rect 32504 15166 32852 15172
rect 32504 15102 32782 15166
rect 32846 15102 32852 15166
rect 32504 15096 32852 15102
rect 32912 15166 34756 15172
rect 32912 15102 34686 15166
rect 34750 15102 34756 15166
rect 32912 15096 34756 15102
rect 39304 15166 39924 15172
rect 39304 15102 39854 15166
rect 39918 15102 39924 15166
rect 39304 15096 39924 15102
rect 28288 15036 28364 15096
rect 28832 15036 28908 15096
rect 28288 14960 28908 15036
rect 30736 15036 30812 15096
rect 31144 15036 31220 15096
rect 30736 14960 31220 15036
rect 31416 15036 31492 15096
rect 32504 15036 32580 15096
rect 31416 14960 32580 15036
rect 39304 15036 39516 15096
rect 39984 15036 40196 15172
rect 39304 14960 40196 15036
rect 25160 14900 25236 14960
rect 25160 14764 25372 14900
rect 34680 14894 34892 14900
rect 34680 14830 34686 14894
rect 34750 14830 34892 14894
rect 15368 14758 15580 14764
rect 15368 14694 15374 14758
rect 15438 14694 15580 14758
rect 15368 14628 15580 14694
rect 16184 14628 16396 14764
rect 17136 14628 17484 14764
rect 17816 14628 18028 14764
rect 18224 14758 19660 14764
rect 18224 14694 19590 14758
rect 19654 14694 19660 14758
rect 18224 14688 19660 14694
rect 25160 14758 25780 14764
rect 25160 14694 25166 14758
rect 25230 14694 25780 14758
rect 25160 14688 25780 14694
rect 34680 14758 34892 14830
rect 39304 14824 39516 14960
rect 39984 14894 40196 14960
rect 39984 14830 40126 14894
rect 40190 14830 40196 14894
rect 39984 14824 40196 14830
rect 34680 14694 34686 14758
rect 34750 14694 34892 14758
rect 34680 14688 34892 14694
rect 15368 14622 17756 14628
rect 15368 14558 17686 14622
rect 17750 14558 17756 14622
rect 15368 14552 17756 14558
rect 17816 14622 18300 14628
rect 17816 14558 18230 14622
rect 18294 14558 18300 14622
rect 17816 14552 18300 14558
rect 25568 14552 25780 14688
rect 34080 14551 34164 14555
rect 34047 14546 34164 14551
rect 34047 14490 34052 14546
rect 34108 14490 34164 14546
rect 34047 14485 34164 14490
rect 34080 14481 34164 14485
rect 17718 14350 19116 14356
rect 17680 14286 17686 14350
rect 17750 14286 19116 14350
rect 17718 14280 19116 14286
rect 18904 14220 19116 14280
rect 19448 14220 19796 14356
rect 20128 14220 20340 14356
rect 20808 14220 21020 14356
rect 21352 14220 21564 14356
rect 18904 14214 21564 14220
rect 18904 14150 19046 14214
rect 19110 14150 20814 14214
rect 20878 14150 21494 14214
rect 21558 14150 21564 14214
rect 18904 14144 21564 14150
rect 22032 14280 22924 14356
rect 22032 14214 22244 14280
rect 22032 14150 22038 14214
rect 22102 14150 22244 14214
rect 22032 14144 22244 14150
rect 22576 14220 22924 14280
rect 23256 14220 23468 14356
rect 23936 14220 24148 14356
rect 24480 14220 24692 14356
rect 35088 14290 35300 14356
rect 35088 14234 35134 14290
rect 35190 14234 35300 14290
rect 22576 14214 23196 14220
rect 22576 14150 22718 14214
rect 22782 14150 23126 14214
rect 23190 14150 23196 14214
rect 22576 14144 23196 14150
rect 23256 14214 23876 14220
rect 23256 14150 23262 14214
rect 23326 14150 23806 14214
rect 23870 14150 23876 14214
rect 23256 14144 23876 14150
rect 23936 14214 24692 14220
rect 23936 14150 23942 14214
rect 24006 14150 24692 14214
rect 33846 14221 33912 14224
rect 34184 14221 34250 14224
rect 33846 14219 34250 14221
rect 33846 14163 33851 14219
rect 33907 14163 34189 14219
rect 34245 14163 34250 14219
rect 33846 14161 34250 14163
rect 33846 14158 33912 14161
rect 34184 14158 34250 14161
rect 35088 14220 35300 14234
rect 23936 14144 24692 14150
rect 35088 14144 43460 14220
rect 1632 13884 1844 13948
rect 1632 13828 1730 13884
rect 1786 13828 1844 13884
rect 1632 13812 1844 13828
rect 3264 13812 3476 14084
rect 3944 13812 4292 14084
rect 1224 13806 4292 13812
rect 1224 13742 1230 13806
rect 1294 13742 4292 13806
rect 1224 13736 4292 13742
rect 9384 14078 10548 14084
rect 9384 14014 10478 14078
rect 10542 14014 10548 14078
rect 9384 14008 10548 14014
rect 9384 13806 9596 14008
rect 41616 13884 41828 13948
rect 41616 13828 41712 13884
rect 41768 13828 41828 13884
rect 41616 13812 41828 13828
rect 9384 13742 9526 13806
rect 9590 13742 9596 13806
rect 9384 13736 9596 13742
rect 19040 13806 19252 13812
rect 19040 13742 19046 13806
rect 19110 13742 19252 13806
rect 19040 13676 19252 13742
rect 19448 13676 19660 13812
rect 19040 13600 19660 13676
rect 20264 13676 20476 13812
rect 20672 13806 20884 13812
rect 20672 13742 20814 13806
rect 20878 13742 20884 13806
rect 20672 13676 20884 13742
rect 20264 13600 20884 13676
rect 21488 13806 22108 13812
rect 21488 13742 21494 13806
rect 21558 13742 22038 13806
rect 22102 13742 22108 13806
rect 21488 13736 22108 13742
rect 21488 13600 21700 13736
rect 21896 13676 22108 13736
rect 22712 13806 22924 13812
rect 22712 13742 22718 13806
rect 22782 13742 22924 13806
rect 21896 13670 22652 13676
rect 21896 13606 22582 13670
rect 22646 13606 22652 13670
rect 21896 13600 22652 13606
rect 22712 13600 22924 13742
rect 23120 13806 23332 13812
rect 23838 13806 24284 13812
rect 23120 13742 23126 13806
rect 23190 13742 23262 13806
rect 23326 13742 23332 13806
rect 23800 13742 23806 13806
rect 23870 13742 23942 13806
rect 24006 13742 24284 13806
rect 23120 13600 23332 13742
rect 23838 13736 24284 13742
rect 23936 13600 24284 13736
rect 41616 13806 42236 13812
rect 41616 13742 42166 13806
rect 42230 13742 42236 13806
rect 41616 13736 42236 13742
rect 41616 13676 41692 13736
rect 39304 13540 39516 13676
rect 39984 13600 41692 13676
rect 39984 13540 40196 13600
rect 32814 13534 34892 13540
rect 32776 13470 32782 13534
rect 32846 13470 34892 13534
rect 32814 13464 34892 13470
rect 39304 13464 40196 13540
rect 34680 13398 34892 13464
rect 34680 13334 34822 13398
rect 34886 13334 34892 13398
rect 34680 13328 34892 13334
rect 9493 13235 9559 13238
rect 15643 13235 15709 13238
rect 9493 13233 15709 13235
rect 9493 13177 9498 13233
rect 9554 13177 15648 13233
rect 15704 13177 15709 13233
rect 9493 13175 15709 13177
rect 9493 13172 9559 13175
rect 15643 13172 15709 13175
rect 2635 12874 2641 12938
rect 2705 12936 2711 12938
rect 2705 12876 19227 12936
rect 2705 12874 2711 12876
rect 40792 12863 40858 12864
rect 40750 12799 40793 12863
rect 40857 12799 40900 12863
rect 40792 12798 40858 12799
rect 33766 12663 33832 12666
rect 34184 12663 34250 12666
rect 33766 12661 34250 12663
rect 19709 12588 19807 12613
rect 20055 12588 20153 12613
rect 20957 12588 21055 12613
rect 21303 12588 21401 12613
rect 22205 12588 22303 12613
rect 22551 12588 22649 12613
rect 23453 12588 23551 12613
rect 23799 12588 23897 12613
rect 33766 12605 33771 12661
rect 33827 12605 34189 12661
rect 34245 12605 34250 12661
rect 33766 12603 34250 12605
rect 33766 12600 33832 12603
rect 34184 12600 34250 12603
rect 35088 12648 43460 12724
rect 35088 12590 35300 12648
rect 3264 12582 3476 12588
rect 3264 12518 3406 12582
rect 3470 12518 3476 12582
rect 3264 12452 3476 12518
rect 3944 12452 4292 12588
rect 3264 12446 4292 12452
rect 3264 12382 4086 12446
rect 4150 12382 4292 12446
rect 3264 12376 4292 12382
rect 9384 12582 10956 12588
rect 9384 12518 10886 12582
rect 10950 12518 10956 12582
rect 9384 12512 10956 12518
rect 19584 12582 25236 12588
rect 19584 12518 19590 12582
rect 19654 12518 20134 12582
rect 20198 12518 25166 12582
rect 25230 12518 25236 12582
rect 19584 12512 25236 12518
rect 35088 12534 35134 12590
rect 35190 12534 35300 12590
rect 35088 12512 35300 12534
rect 9384 12446 9596 12512
rect 9384 12382 9390 12446
rect 9454 12382 9596 12446
rect 9384 12376 9596 12382
rect 1224 12310 1844 12316
rect 1224 12246 1230 12310
rect 1294 12246 1844 12310
rect 1224 12240 1844 12246
rect 1632 12204 1844 12240
rect 1632 12148 1730 12204
rect 1786 12148 1844 12204
rect 39304 12180 39516 12316
rect 39984 12310 40196 12316
rect 39984 12246 40126 12310
rect 40190 12246 40196 12310
rect 39984 12180 40196 12246
rect 1632 12104 1844 12148
rect 34680 12174 34892 12180
rect 34680 12110 34686 12174
rect 34750 12110 34892 12174
rect 19584 11772 19796 11908
rect 20128 11832 21564 11908
rect 20128 11772 20340 11832
rect 19584 11766 20340 11772
rect 19584 11702 20270 11766
rect 20334 11702 20340 11766
rect 19584 11696 20340 11702
rect 20808 11696 21020 11832
rect 21352 11772 21564 11832
rect 22032 11772 22244 11908
rect 22576 11902 23604 11908
rect 22576 11838 22582 11902
rect 22646 11838 23604 11902
rect 22576 11832 23604 11838
rect 22576 11772 22788 11832
rect 21352 11696 22788 11772
rect 23256 11772 23604 11832
rect 23800 11772 24012 11908
rect 34680 11902 34892 12110
rect 39304 12104 40196 12180
rect 41616 12310 42236 12316
rect 41616 12246 42166 12310
rect 42230 12246 42236 12310
rect 41616 12240 42236 12246
rect 41616 12204 41828 12240
rect 41616 12148 41712 12204
rect 41768 12148 41828 12204
rect 41616 12104 41828 12148
rect 34680 11838 34686 11902
rect 34750 11838 34892 11902
rect 34680 11832 34892 11838
rect 23256 11696 24012 11772
rect 35088 11462 35300 11500
rect 35088 11406 35134 11462
rect 35190 11406 35300 11462
rect 33686 11393 33752 11396
rect 34184 11393 34250 11396
rect 33686 11391 34250 11393
rect 33686 11335 33691 11391
rect 33747 11335 34189 11391
rect 34245 11335 34250 11391
rect 33686 11333 34250 11335
rect 33686 11330 33752 11333
rect 34184 11330 34250 11333
rect 35088 11364 35300 11406
rect 35088 11288 43460 11364
rect 3264 11152 4292 11228
rect 3264 11086 3476 11152
rect 3264 11022 3270 11086
rect 3334 11022 3476 11086
rect 3264 11016 3476 11022
rect 3944 11016 4292 11152
rect 9384 11222 9596 11228
rect 9384 11158 9526 11222
rect 9590 11158 9596 11222
rect 9384 11086 9596 11158
rect 9384 11022 9526 11086
rect 9590 11022 9596 11086
rect 9384 11016 9596 11022
rect 19584 11086 24012 11092
rect 19584 11022 20270 11086
rect 20334 11022 24012 11086
rect 19584 11016 24012 11022
rect 19639 10903 19737 11016
rect 19992 10950 20223 11016
rect 19992 10886 19998 10950
rect 20062 10903 20223 10950
rect 20887 10903 20985 11016
rect 20062 10886 20204 10903
rect 19992 10880 20204 10886
rect 21352 10880 21564 11016
rect 22135 10903 22233 11016
rect 22621 10903 22788 11016
rect 23383 10903 23481 11016
rect 23869 10903 24012 11016
rect 22712 10880 22788 10903
rect 23936 10880 24012 10903
rect 19312 10814 19796 10820
rect 19312 10750 19726 10814
rect 19790 10750 19796 10814
rect 19312 10744 19796 10750
rect 20264 10744 20476 10820
rect 20536 10814 21020 10820
rect 20536 10750 20950 10814
rect 21014 10750 21020 10814
rect 20536 10744 21020 10750
rect 19312 10677 19524 10744
rect 20400 10698 20476 10744
rect 19992 10679 20204 10684
rect 19312 10621 19406 10677
rect 19462 10621 19524 10677
rect 1632 10542 3340 10548
rect 1632 10524 3270 10542
rect 1632 10468 1730 10524
rect 1786 10478 3270 10524
rect 3334 10478 3340 10542
rect 1786 10472 3340 10478
rect 19312 10472 19524 10621
rect 19639 10548 19737 10679
rect 19992 10678 20223 10679
rect 19992 10614 20134 10678
rect 20198 10614 20223 10678
rect 19992 10581 20223 10614
rect 20379 10677 20477 10698
rect 20633 10684 20748 10744
rect 21624 10698 21700 10820
rect 21896 10814 22516 10820
rect 21896 10750 22446 10814
rect 22510 10750 22516 10814
rect 21896 10744 22516 10750
rect 21896 10698 21972 10744
rect 20379 10621 20400 10677
rect 20456 10621 20477 10677
rect 20379 10600 20477 10621
rect 20536 10677 20748 10684
rect 20536 10621 20654 10677
rect 20710 10621 20748 10677
rect 20536 10608 20748 10621
rect 19992 10548 20204 10581
rect 20400 10548 20476 10600
rect 20633 10548 20748 10608
rect 19639 10542 20204 10548
rect 19639 10510 20134 10542
rect 19720 10478 20134 10510
rect 20198 10478 20204 10542
rect 19720 10472 20204 10478
rect 20264 10542 20476 10548
rect 20264 10478 20270 10542
rect 20334 10478 20476 10542
rect 20264 10472 20476 10478
rect 20536 10472 20748 10548
rect 20887 10548 20985 10679
rect 21352 10548 21564 10684
rect 20887 10542 21564 10548
rect 20887 10510 21494 10542
rect 20944 10478 21494 10510
rect 21558 10478 21564 10542
rect 20944 10472 21564 10478
rect 21624 10677 21725 10698
rect 21624 10621 21648 10677
rect 21704 10621 21725 10677
rect 21624 10600 21725 10621
rect 21881 10677 21979 10698
rect 22712 10679 22788 10684
rect 21881 10621 21902 10677
rect 21958 10621 21979 10677
rect 21881 10600 21979 10621
rect 21624 10542 21700 10600
rect 21624 10478 21630 10542
rect 21694 10478 21700 10542
rect 21624 10472 21700 10478
rect 21896 10472 21972 10600
rect 22135 10548 22233 10679
rect 22621 10548 22788 10679
rect 22135 10542 22788 10548
rect 22135 10510 22174 10542
rect 22168 10478 22174 10510
rect 22238 10478 22718 10542
rect 22782 10478 22788 10542
rect 22168 10472 22788 10478
rect 22848 10677 23060 10820
rect 22848 10621 22896 10677
rect 22952 10621 23060 10677
rect 22848 10542 23060 10621
rect 22848 10478 22854 10542
rect 22918 10478 23060 10542
rect 22848 10472 23060 10478
rect 23120 10814 23740 10820
rect 23120 10750 23670 10814
rect 23734 10750 23740 10814
rect 23120 10744 23740 10750
rect 23120 10677 23227 10744
rect 23936 10679 24012 10684
rect 23120 10621 23150 10677
rect 23206 10621 23227 10677
rect 23120 10600 23227 10621
rect 23120 10472 23196 10600
rect 23383 10548 23481 10679
rect 23869 10548 24012 10679
rect 23383 10542 24012 10548
rect 23383 10510 23398 10542
rect 23392 10478 23398 10510
rect 23462 10478 23942 10542
rect 24006 10478 24012 10542
rect 23392 10472 24012 10478
rect 24072 10677 24284 10820
rect 24072 10621 24144 10677
rect 24200 10621 24284 10677
rect 24072 10542 24284 10621
rect 24072 10478 24078 10542
rect 24142 10478 24284 10542
rect 24072 10472 24284 10478
rect 34680 10678 34892 10684
rect 34680 10614 34822 10678
rect 34886 10614 34892 10678
rect 34680 10472 34892 10614
rect 41616 10524 41828 10548
rect 1786 10468 1844 10472
rect 1632 10412 1844 10468
rect 1224 10406 1844 10412
rect 1224 10342 1230 10406
rect 1294 10342 1844 10406
rect 9493 10444 9559 10447
rect 17294 10444 17360 10447
rect 9493 10442 17360 10444
rect 9493 10386 9498 10442
rect 9554 10386 17299 10442
rect 17355 10386 17360 10442
rect 9493 10384 17360 10386
rect 9493 10381 9559 10384
rect 17294 10381 17360 10384
rect 1224 10336 1844 10342
rect 22712 10276 22788 10472
rect 41616 10468 41712 10524
rect 41768 10468 41828 10524
rect 41616 10412 41828 10468
rect 41616 10406 42236 10412
rect 41616 10342 42166 10406
rect 42230 10342 42236 10406
rect 41616 10336 42236 10342
rect 22712 10270 23468 10276
rect 22712 10206 23398 10270
rect 23462 10206 23468 10270
rect 22712 10200 23468 10206
rect 21526 10134 21972 10140
rect 21488 10070 21494 10134
rect 21558 10070 21972 10134
rect 21526 10064 21972 10070
rect 21896 10004 21972 10064
rect 19448 9998 20340 10004
rect 19448 9934 20134 9998
rect 20198 9934 20340 9998
rect 19448 9928 20340 9934
rect 3264 9726 4292 9732
rect 3264 9662 4086 9726
rect 4150 9662 4292 9726
rect 3264 9656 4292 9662
rect 3264 9520 3476 9656
rect 3944 9520 4292 9656
rect 9384 9726 9596 9732
rect 9384 9662 9390 9726
rect 9454 9662 9596 9726
rect 9384 9590 9596 9662
rect 19448 9656 19660 9928
rect 19992 9726 20340 9928
rect 19992 9662 20134 9726
rect 20198 9662 20340 9726
rect 19992 9656 20340 9662
rect 20672 9726 20884 10004
rect 20672 9662 20814 9726
rect 20878 9662 20884 9726
rect 20672 9656 20884 9662
rect 21352 9868 21564 10004
rect 21896 9998 22244 10004
rect 21896 9934 22174 9998
rect 22238 9934 22244 9998
rect 21896 9868 22244 9934
rect 21352 9792 22244 9868
rect 21352 9656 21564 9792
rect 21896 9656 22244 9792
rect 22576 9998 22788 10004
rect 22576 9934 22718 9998
rect 22782 9934 22788 9998
rect 22576 9656 22788 9934
rect 23256 9732 23468 10004
rect 23800 9998 24012 10004
rect 23800 9934 23942 9998
rect 24006 9934 24012 9998
rect 23800 9732 24012 9934
rect 33606 9835 33672 9838
rect 34184 9835 34250 9838
rect 33606 9833 34250 9835
rect 33606 9777 33611 9833
rect 33667 9777 34189 9833
rect 34245 9777 34250 9833
rect 33606 9775 34250 9777
rect 33606 9772 33672 9775
rect 34184 9772 34250 9775
rect 23256 9726 24012 9732
rect 23256 9662 23262 9726
rect 23326 9662 24012 9726
rect 23256 9656 24012 9662
rect 35088 9762 35300 9868
rect 35088 9706 35134 9762
rect 35190 9732 35300 9762
rect 35190 9706 43460 9732
rect 35088 9656 43460 9706
rect 9384 9526 9390 9590
rect 9454 9526 9596 9590
rect 9384 9520 9596 9526
rect 19856 9590 20068 9596
rect 19856 9526 19998 9590
rect 20062 9526 20068 9590
rect 19856 9520 20068 9526
rect 19856 9460 19932 9520
rect 19448 9384 19932 9460
rect 19448 9324 19660 9384
rect 19992 9324 20340 9460
rect 20672 9384 21564 9460
rect 20672 9324 20884 9384
rect 19448 9318 20884 9324
rect 19448 9254 20678 9318
rect 20742 9254 20884 9318
rect 19448 9248 20884 9254
rect 21352 9324 21564 9384
rect 21896 9324 22244 9460
rect 22576 9324 22788 9460
rect 23256 9324 23468 9460
rect 23800 9324 24012 9460
rect 21352 9248 24012 9324
rect 34680 9318 34892 9324
rect 34680 9254 34686 9318
rect 34750 9254 34892 9318
rect 19584 9052 19796 9188
rect 19992 9182 20204 9188
rect 19992 9118 20134 9182
rect 20198 9118 20204 9182
rect 19992 9052 20204 9118
rect 9493 8993 9559 8996
rect 17542 8993 17608 8996
rect 9493 8991 17608 8993
rect 9493 8935 9498 8991
rect 9554 8935 17547 8991
rect 17603 8935 17608 8991
rect 9493 8933 17608 8935
rect 9493 8930 9559 8933
rect 17542 8930 17608 8933
rect 19584 8976 20204 9052
rect 20808 9182 21020 9188
rect 20808 9118 20814 9182
rect 20878 9118 21020 9182
rect 20808 9052 21020 9118
rect 21216 9052 21428 9188
rect 20808 8976 21428 9052
rect 22032 9112 22652 9188
rect 22032 8976 22244 9112
rect 22440 8976 22652 9112
rect 23256 9182 23604 9188
rect 23256 9118 23262 9182
rect 23326 9118 23604 9182
rect 23256 9052 23604 9118
rect 23664 9052 23876 9188
rect 34680 9112 34892 9254
rect 19584 8916 19660 8976
rect 1224 8910 1844 8916
rect 1224 8846 1230 8910
rect 1294 8846 1844 8910
rect 1224 8844 1844 8846
rect 1224 8840 1730 8844
rect 1632 8788 1730 8840
rect 1786 8788 1844 8844
rect 1632 8780 1844 8788
rect 19448 8780 19660 8916
rect 1632 8774 3340 8780
rect 19078 8774 19660 8780
rect 1632 8710 3270 8774
rect 3334 8710 3340 8774
rect 19040 8710 19046 8774
rect 19110 8710 19660 8774
rect 1632 8704 3340 8710
rect 19078 8704 19660 8710
rect 19992 8916 20068 8976
rect 20808 8916 20884 8976
rect 19992 8840 20884 8916
rect 19992 8704 20340 8840
rect 20672 8704 20884 8840
rect 21352 8916 21428 8976
rect 22168 8916 22244 8976
rect 21352 8780 21564 8916
rect 21896 8780 22244 8916
rect 21352 8704 22244 8780
rect 22576 8916 22652 8976
rect 23120 8976 23876 9052
rect 23120 8916 23196 8976
rect 22576 8840 23196 8916
rect 23256 8916 23332 8976
rect 23800 8916 23876 8976
rect 22576 8704 22788 8840
rect 23256 8704 23468 8916
rect 23800 8780 24012 8916
rect 41616 8844 41828 8916
rect 41616 8788 41712 8844
rect 41768 8788 41828 8844
rect 41616 8780 41828 8788
rect 23800 8774 24556 8780
rect 23800 8710 24486 8774
rect 24550 8710 24556 8774
rect 23800 8704 24556 8710
rect 41616 8774 42236 8780
rect 41616 8710 42166 8774
rect 42230 8710 42236 8774
rect 41616 8704 42236 8710
rect 19350 8502 24420 8508
rect 19312 8438 19318 8502
rect 19382 8438 20678 8502
rect 20742 8438 24350 8502
rect 24414 8438 24420 8502
rect 19350 8432 24420 8438
rect 19534 8401 19632 8432
rect 20106 8401 20204 8432
rect 20782 8401 20880 8432
rect 21354 8401 21452 8432
rect 22030 8401 22128 8432
rect 22602 8401 22700 8432
rect 23278 8401 23376 8432
rect 23850 8401 23948 8432
rect 3264 8366 3476 8372
rect 3264 8302 3270 8366
rect 3334 8302 3476 8366
rect 3264 8236 3476 8302
rect 3944 8236 4292 8372
rect 3264 8160 4292 8236
rect 9384 8366 9596 8372
rect 9384 8302 9526 8366
rect 9590 8302 9596 8366
rect 9384 8230 9596 8302
rect 9384 8166 9526 8230
rect 9590 8166 9596 8230
rect 9384 8160 9596 8166
rect 17816 8094 19388 8100
rect 17816 8030 19318 8094
rect 19382 8030 19388 8094
rect 17816 8024 19388 8030
rect 24208 8094 24420 8100
rect 24208 8030 24350 8094
rect 24414 8030 24420 8094
rect 17816 7888 18028 8024
rect 24208 7888 24420 8030
rect 9493 7595 9559 7598
rect 17418 7595 17484 7598
rect 9493 7593 17484 7595
rect 9493 7537 9498 7593
rect 9554 7537 17423 7593
rect 17479 7537 17484 7593
rect 9493 7535 17484 7537
rect 9493 7532 9559 7535
rect 17418 7532 17484 7535
rect 1632 7164 1844 7284
rect 1632 7148 1730 7164
rect 1224 7142 1730 7148
rect 1224 7078 1230 7142
rect 1294 7108 1730 7142
rect 1786 7108 1844 7164
rect 1294 7078 1844 7108
rect 1224 7072 1844 7078
rect 41616 7164 41828 7284
rect 41616 7108 41712 7164
rect 41768 7148 41828 7164
rect 41768 7142 42236 7148
rect 41768 7108 42166 7142
rect 41616 7078 42166 7108
rect 42230 7078 42236 7142
rect 41616 7072 42236 7078
rect 9384 7006 9596 7012
rect 9384 6942 9390 7006
rect 9454 6942 9596 7006
rect 9384 6734 9596 6942
rect 17816 7006 19116 7012
rect 17816 6942 19046 7006
rect 19110 6942 19116 7006
rect 17816 6936 19116 6942
rect 24208 7006 24518 7012
rect 24208 6942 24486 7006
rect 24550 6942 24556 7006
rect 24208 6936 24518 6942
rect 17816 6800 18028 6936
rect 24208 6800 24420 6936
rect 9384 6670 9526 6734
rect 9590 6670 9596 6734
rect 9384 6664 9596 6670
rect 544 5646 1980 5652
rect 544 5582 550 5646
rect 614 5582 1980 5646
rect 544 5576 1980 5582
rect 1904 5516 1980 5576
rect 1632 5484 1844 5516
rect 1632 5428 1730 5484
rect 1786 5428 1844 5484
rect 1904 5440 2796 5516
rect 1632 5380 1844 5428
rect 1224 5374 1844 5380
rect 1224 5310 1230 5374
rect 1294 5310 1844 5374
rect 1224 5304 1844 5310
rect 2584 5304 2796 5440
rect 9384 5510 9596 5516
rect 9384 5446 9390 5510
rect 9454 5446 9596 5510
rect 9384 5380 9596 5446
rect 9248 5374 9596 5380
rect 9248 5310 9254 5374
rect 9318 5310 9596 5374
rect 9248 5304 9596 5310
rect 41616 5484 41828 5516
rect 41616 5428 41712 5484
rect 41768 5428 41828 5484
rect 41616 5380 41828 5428
rect 41616 5374 42236 5380
rect 41616 5310 42166 5374
rect 42230 5310 42236 5374
rect 41616 5304 42236 5310
rect 2720 4892 3068 4972
rect 2720 4836 2858 4892
rect 2914 4836 3068 4892
rect 0 4760 3068 4836
rect 2584 3944 2796 4156
rect 9384 4150 9596 4156
rect 9384 4086 9526 4150
rect 9590 4086 9596 4150
rect 9384 4020 9596 4086
rect 11152 4080 12588 4156
rect 11152 4020 11364 4080
rect 9384 4014 11364 4020
rect 9384 3950 9390 4014
rect 9454 3950 11364 4014
rect 9384 3944 11364 3950
rect 12376 4020 12588 4080
rect 13464 4080 17212 4156
rect 13464 4020 13676 4080
rect 12376 3944 13676 4020
rect 14688 3944 14900 4080
rect 15776 3944 16124 4080
rect 17000 4020 17212 4080
rect 18224 4080 19524 4156
rect 18224 4020 18436 4080
rect 17000 3944 18436 4020
rect 19312 4020 19524 4080
rect 20536 4080 24284 4156
rect 20536 4020 20748 4080
rect 19312 3944 20748 4020
rect 21624 3944 21972 4080
rect 22848 3944 23060 4080
rect 24072 3944 24284 4080
rect 2584 3884 2660 3944
rect 1224 3878 2660 3884
rect 1224 3814 1230 3878
rect 1294 3814 2660 3878
rect 1224 3808 2660 3814
rect 41616 3878 42236 3884
rect 41616 3814 42166 3878
rect 42230 3814 42236 3878
rect 41616 3808 42236 3814
rect 1632 3804 1844 3808
rect 1632 3748 1730 3804
rect 1786 3748 1844 3804
rect 1632 3672 1844 3748
rect 41616 3804 41828 3808
rect 41616 3748 41712 3804
rect 41768 3748 41828 3804
rect 41616 3672 41828 3748
rect 2720 3192 3068 3340
rect 2720 3136 2858 3192
rect 2914 3136 3068 3192
rect 2720 3068 3068 3136
rect 5984 3297 6196 3340
rect 5984 3241 6079 3297
rect 6135 3241 6196 3297
rect 5984 3198 6196 3241
rect 5984 3134 5990 3198
rect 6054 3134 6196 3198
rect 5984 3128 6196 3134
rect 10744 3198 10956 3340
rect 10744 3134 10750 3198
rect 10814 3192 10956 3198
rect 10814 3136 10836 3192
rect 10892 3136 10956 3192
rect 10814 3134 10956 3136
rect 10744 3128 10956 3134
rect 11968 3198 12180 3340
rect 13192 3213 13268 3340
rect 14416 3213 14492 3340
rect 15504 3213 15716 3340
rect 16728 3213 16804 3340
rect 11968 3192 12110 3198
rect 11968 3136 12004 3192
rect 12060 3136 12110 3192
rect 11968 3134 12110 3136
rect 12174 3134 12180 3198
rect 11968 3128 12180 3134
rect 13151 3198 13268 3213
rect 13151 3192 13198 3198
rect 13151 3136 13172 3192
rect 13151 3134 13198 3136
rect 13262 3134 13268 3198
rect 13151 3128 13268 3134
rect 14319 3198 14492 3213
rect 14319 3192 14422 3198
rect 14319 3136 14340 3192
rect 14396 3136 14422 3192
rect 14319 3134 14422 3136
rect 14486 3134 14492 3198
rect 14319 3128 14492 3134
rect 15487 3198 15716 3213
rect 15487 3192 15510 3198
rect 15487 3136 15508 3192
rect 15487 3134 15510 3136
rect 15574 3134 15716 3198
rect 15487 3128 15716 3134
rect 16655 3198 16804 3213
rect 16655 3192 16734 3198
rect 16655 3136 16676 3192
rect 16732 3136 16734 3192
rect 16655 3134 16734 3136
rect 16798 3134 16804 3198
rect 16655 3128 16804 3134
rect 17816 3198 18028 3340
rect 19040 3213 19116 3340
rect 17816 3192 17958 3198
rect 17816 3136 17844 3192
rect 17900 3136 17958 3192
rect 17816 3134 17958 3136
rect 18022 3134 18028 3198
rect 17816 3128 18028 3134
rect 18991 3198 19116 3213
rect 18991 3192 19046 3198
rect 18991 3136 19012 3192
rect 18991 3134 19046 3136
rect 19110 3134 19116 3198
rect 18991 3128 19116 3134
rect 20128 3198 20340 3340
rect 21352 3213 21428 3340
rect 22576 3213 22652 3340
rect 23664 3213 23876 3340
rect 20128 3192 20270 3198
rect 20128 3136 20180 3192
rect 20236 3136 20270 3192
rect 20128 3134 20270 3136
rect 20334 3134 20340 3198
rect 20128 3128 20340 3134
rect 21327 3198 21428 3213
rect 21327 3192 21358 3198
rect 21327 3136 21348 3192
rect 21327 3134 21358 3136
rect 21422 3134 21428 3198
rect 21327 3128 21428 3134
rect 22495 3198 22652 3213
rect 22495 3192 22582 3198
rect 22495 3136 22516 3192
rect 22572 3136 22582 3192
rect 22495 3134 22582 3136
rect 22646 3134 22652 3198
rect 22495 3128 22652 3134
rect 23663 3198 23876 3213
rect 23663 3192 23806 3198
rect 23663 3136 23684 3192
rect 23740 3136 23806 3192
rect 23663 3134 23806 3136
rect 23870 3134 23876 3198
rect 23663 3128 23876 3134
rect 10815 3115 10913 3128
rect 11983 3115 12081 3128
rect 13151 3115 13249 3128
rect 14319 3115 14417 3128
rect 15487 3115 15585 3128
rect 16655 3115 16753 3128
rect 17823 3115 17921 3128
rect 18991 3115 19089 3128
rect 20159 3115 20257 3128
rect 21327 3115 21425 3128
rect 22495 3115 22593 3128
rect 23663 3115 23761 3128
rect 0 2992 3068 3068
rect 9577 2938 9643 2941
rect 9577 2936 20038 2938
rect 9577 2880 9582 2936
rect 9638 2880 20038 2936
rect 9577 2878 20038 2880
rect 9577 2875 9643 2878
rect 2584 2524 2796 2660
rect 9286 2654 9596 2660
rect 9248 2590 9254 2654
rect 9318 2590 9596 2654
rect 9286 2584 9596 2590
rect 544 2518 2796 2524
rect 544 2454 550 2518
rect 614 2454 2796 2518
rect 544 2448 2796 2454
rect 9384 2524 9596 2584
rect 11152 2584 13676 2660
rect 11152 2524 11364 2584
rect 9384 2518 11364 2524
rect 9384 2454 9526 2518
rect 9590 2454 11364 2518
rect 9384 2448 11364 2454
rect 12376 2448 12588 2584
rect 13464 2524 13676 2584
rect 14688 2584 17212 2660
rect 14688 2524 14900 2584
rect 13464 2448 14900 2524
rect 15776 2448 16124 2584
rect 17000 2524 17212 2584
rect 18224 2584 19524 2660
rect 18224 2524 18436 2584
rect 17000 2448 18436 2524
rect 19312 2524 19524 2584
rect 20536 2584 21972 2660
rect 20536 2524 20748 2584
rect 19312 2448 20748 2524
rect 21624 2524 21972 2584
rect 22848 2584 24284 2660
rect 22848 2524 23060 2584
rect 21624 2448 23060 2524
rect 24072 2448 24284 2584
rect 1632 2124 1844 2252
rect 1632 2068 1730 2124
rect 1786 2116 1844 2124
rect 41616 2124 41828 2252
rect 1786 2110 2116 2116
rect 1786 2068 2046 2110
rect 1632 2046 2046 2068
rect 2110 2046 2116 2110
rect 1632 2040 2116 2046
rect 41616 2068 41712 2124
rect 41768 2116 41828 2124
rect 41768 2110 42236 2116
rect 41768 2068 42166 2110
rect 41616 2046 42166 2068
rect 42230 2046 42236 2110
rect 41616 2040 42236 2046
rect 2040 1838 2252 1844
rect 2040 1774 2046 1838
rect 2110 1788 2252 1838
rect 2040 1732 2066 1774
rect 2122 1732 2252 1788
rect 2040 1702 2252 1732
rect 2040 1638 2182 1702
rect 2246 1638 2252 1702
rect 2040 1632 2252 1638
rect 3672 1788 3884 1844
rect 3672 1732 3746 1788
rect 3802 1732 3884 1788
rect 3672 1702 3884 1732
rect 3672 1638 3814 1702
rect 3878 1638 3884 1702
rect 3672 1632 3884 1638
rect 5304 1788 5516 1844
rect 5304 1732 5426 1788
rect 5482 1732 5516 1788
rect 5304 1702 5516 1732
rect 5304 1638 5446 1702
rect 5510 1638 5516 1702
rect 5304 1632 5516 1638
rect 7072 1788 7284 1844
rect 7072 1732 7106 1788
rect 7162 1732 7284 1788
rect 7072 1702 7284 1732
rect 7072 1638 7078 1702
rect 7142 1638 7284 1702
rect 7072 1632 7284 1638
rect 8704 1838 9460 1844
rect 8704 1788 9390 1838
rect 8704 1732 8786 1788
rect 8842 1774 9390 1788
rect 9454 1774 9460 1838
rect 8842 1768 9460 1774
rect 10336 1788 10548 1844
rect 8842 1732 8916 1768
rect 8704 1702 8916 1732
rect 8704 1638 8710 1702
rect 8774 1638 8916 1702
rect 8704 1632 8916 1638
rect 10336 1732 10466 1788
rect 10522 1732 10548 1788
rect 10336 1702 10548 1732
rect 10336 1638 10342 1702
rect 10406 1638 10548 1702
rect 10336 1632 10548 1638
rect 12104 1788 12316 1844
rect 12104 1732 12146 1788
rect 12202 1732 12316 1788
rect 12104 1702 12316 1732
rect 12104 1638 12246 1702
rect 12310 1638 12316 1702
rect 12104 1632 12316 1638
rect 13736 1788 13948 1844
rect 13736 1732 13826 1788
rect 13882 1732 13948 1788
rect 13736 1702 13948 1732
rect 13736 1638 13742 1702
rect 13806 1638 13948 1702
rect 13736 1632 13948 1638
rect 15368 1788 15716 1844
rect 15368 1732 15506 1788
rect 15562 1732 15716 1788
rect 15368 1702 15716 1732
rect 15368 1638 15374 1702
rect 15438 1638 15716 1702
rect 15368 1632 15716 1638
rect 17136 1788 17348 1844
rect 17136 1732 17186 1788
rect 17242 1732 17348 1788
rect 17136 1702 17348 1732
rect 17136 1638 17278 1702
rect 17342 1638 17348 1702
rect 17136 1632 17348 1638
rect 18768 1788 18980 1844
rect 18768 1732 18866 1788
rect 18922 1732 18980 1788
rect 18768 1702 18980 1732
rect 18768 1638 18774 1702
rect 18838 1638 18980 1702
rect 18768 1632 18980 1638
rect 20400 1788 20748 1844
rect 20400 1732 20546 1788
rect 20602 1732 20748 1788
rect 20400 1702 20748 1732
rect 20400 1638 20678 1702
rect 20742 1638 20748 1702
rect 20400 1632 20748 1638
rect 22168 1788 22380 1844
rect 22168 1732 22226 1788
rect 22282 1732 22380 1788
rect 22168 1702 22380 1732
rect 23800 1788 24012 1844
rect 23800 1732 23906 1788
rect 23962 1732 24012 1788
rect 23800 1708 24012 1732
rect 22168 1638 22310 1702
rect 22374 1638 22380 1702
rect 22168 1632 22380 1638
rect 23528 1702 24012 1708
rect 23528 1638 23534 1702
rect 23598 1638 24012 1702
rect 23528 1632 24012 1638
rect 25432 1788 25780 1844
rect 25432 1732 25586 1788
rect 25642 1732 25780 1788
rect 25432 1702 25780 1732
rect 25432 1638 25438 1702
rect 25502 1638 25780 1702
rect 25432 1632 25780 1638
rect 27200 1788 27412 1844
rect 27200 1732 27266 1788
rect 27322 1732 27412 1788
rect 27200 1702 27412 1732
rect 27200 1638 27342 1702
rect 27406 1638 27412 1702
rect 27200 1632 27412 1638
rect 28832 1788 29044 1844
rect 28832 1732 28946 1788
rect 29002 1732 29044 1788
rect 28832 1702 29044 1732
rect 28832 1638 28974 1702
rect 29038 1638 29044 1702
rect 28832 1632 29044 1638
rect 30600 1788 30812 1844
rect 30600 1732 30626 1788
rect 30682 1732 30812 1788
rect 30600 1702 30812 1732
rect 30600 1638 30606 1702
rect 30670 1638 30812 1702
rect 30600 1632 30812 1638
rect 32232 1788 32444 1844
rect 32232 1732 32306 1788
rect 32362 1732 32444 1788
rect 32232 1702 32444 1732
rect 32232 1638 32238 1702
rect 32302 1638 32444 1702
rect 32232 1632 32444 1638
rect 33864 1788 34076 1844
rect 33864 1732 33986 1788
rect 34042 1732 34076 1788
rect 33864 1702 34076 1732
rect 33864 1638 34006 1702
rect 34070 1638 34076 1702
rect 33864 1632 34076 1638
rect 35632 1788 35844 1844
rect 35632 1732 35666 1788
rect 35722 1732 35844 1788
rect 35632 1702 35844 1732
rect 35632 1638 35638 1702
rect 35702 1638 35844 1702
rect 35632 1632 35844 1638
rect 37264 1788 37476 1844
rect 37264 1732 37346 1788
rect 37402 1732 37476 1788
rect 37264 1702 37476 1732
rect 37264 1638 37406 1702
rect 37470 1638 37476 1702
rect 37264 1632 37476 1638
rect 38896 1788 39108 1844
rect 38896 1732 39026 1788
rect 39082 1732 39108 1788
rect 38896 1702 39108 1732
rect 38896 1638 39038 1702
rect 39102 1638 39108 1702
rect 38896 1632 39108 1638
rect 40664 1788 40876 1844
rect 40664 1732 40706 1788
rect 40762 1732 40876 1788
rect 40664 1702 40876 1732
rect 40664 1638 40806 1702
rect 40870 1638 40876 1702
rect 40664 1632 40876 1638
rect 952 1294 42508 1300
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 2182 1294
rect 2246 1230 3814 1294
rect 3878 1230 5446 1294
rect 5510 1230 7078 1294
rect 7142 1230 8710 1294
rect 8774 1230 10342 1294
rect 10406 1230 12246 1294
rect 12310 1230 13742 1294
rect 13806 1230 15374 1294
rect 15438 1230 17278 1294
rect 17342 1230 18774 1294
rect 18838 1230 20678 1294
rect 20742 1230 22310 1294
rect 22374 1230 23534 1294
rect 23598 1230 25438 1294
rect 25502 1230 27342 1294
rect 27406 1230 28974 1294
rect 29038 1230 30606 1294
rect 30670 1230 32238 1294
rect 32302 1230 34006 1294
rect 34070 1230 35638 1294
rect 35702 1230 37406 1294
rect 37470 1230 39038 1294
rect 39102 1230 40806 1294
rect 40870 1230 42166 1294
rect 42230 1230 42302 1294
rect 42366 1230 42438 1294
rect 42502 1230 42508 1294
rect 952 1158 42508 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 42166 1158
rect 42230 1094 42302 1158
rect 42366 1094 42438 1158
rect 42502 1094 42508 1158
rect 952 1022 42508 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 42166 1022
rect 42230 958 42302 1022
rect 42366 958 42438 1022
rect 42502 958 42508 1022
rect 952 952 42508 958
rect 272 614 43188 620
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 9526 614
rect 9590 550 42846 614
rect 42910 550 42982 614
rect 43046 550 43118 614
rect 43182 550 43188 614
rect 272 478 43188 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 42846 478
rect 42910 414 42982 478
rect 43046 414 43118 478
rect 43182 414 43188 478
rect 272 342 43188 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 42846 342
rect 42910 278 42982 342
rect 43046 278 43118 342
rect 43182 278 43188 342
rect 272 272 43188 278
<< via3 >>
rect 278 32782 342 32846
rect 414 32782 478 32846
rect 550 32782 614 32846
rect 42846 32782 42910 32846
rect 42982 32782 43046 32846
rect 43118 32782 43182 32846
rect 278 32646 342 32710
rect 414 32646 478 32710
rect 550 32646 614 32710
rect 42846 32646 42910 32710
rect 42982 32646 43046 32710
rect 43118 32646 43182 32710
rect 278 32510 342 32574
rect 414 32510 478 32574
rect 550 32510 614 32574
rect 34278 32510 34342 32574
rect 42846 32510 42910 32574
rect 42982 32510 43046 32574
rect 43118 32510 43182 32574
rect 958 32102 1022 32166
rect 1094 32102 1158 32166
rect 1230 32102 1294 32166
rect 42166 32102 42230 32166
rect 42302 32102 42366 32166
rect 42438 32102 42502 32166
rect 958 31966 1022 32030
rect 1094 31966 1158 32030
rect 1230 31966 1294 32030
rect 42166 31966 42230 32030
rect 42302 31966 42366 32030
rect 42438 31966 42502 32030
rect 958 31830 1022 31894
rect 1094 31830 1158 31894
rect 1230 31830 1294 31894
rect 2182 31830 2246 31894
rect 3814 31830 3878 31894
rect 5310 31830 5374 31894
rect 7078 31830 7142 31894
rect 8710 31830 8774 31894
rect 10342 31830 10406 31894
rect 12110 31830 12174 31894
rect 13742 31830 13806 31894
rect 15646 31830 15710 31894
rect 17278 31830 17342 31894
rect 18774 31830 18838 31894
rect 20270 31830 20334 31894
rect 22310 31830 22374 31894
rect 23806 31830 23870 31894
rect 25574 31830 25638 31894
rect 27206 31830 27270 31894
rect 28974 31830 29038 31894
rect 30606 31830 30670 31894
rect 32238 31830 32302 31894
rect 34006 31830 34070 31894
rect 35638 31830 35702 31894
rect 37270 31830 37334 31894
rect 38902 31830 38966 31894
rect 40670 31830 40734 31894
rect 42166 31830 42230 31894
rect 42302 31830 42366 31894
rect 42438 31830 42502 31894
rect 2182 31422 2246 31486
rect 3814 31422 3878 31486
rect 5310 31422 5374 31486
rect 7078 31422 7142 31486
rect 8710 31422 8774 31486
rect 10342 31422 10406 31486
rect 12110 31422 12174 31486
rect 13742 31422 13806 31486
rect 15646 31422 15710 31486
rect 17278 31422 17342 31486
rect 18774 31422 18838 31486
rect 20270 31422 20334 31486
rect 22310 31422 22374 31486
rect 23806 31422 23870 31486
rect 25574 31422 25638 31486
rect 27206 31422 27270 31486
rect 28974 31422 29038 31486
rect 30606 31422 30670 31486
rect 32238 31422 32302 31486
rect 34006 31422 34070 31486
rect 35638 31422 35702 31486
rect 34142 31286 34206 31350
rect 37270 31422 37334 31486
rect 38902 31422 38966 31486
rect 40670 31422 40734 31486
rect 1230 30742 1294 30806
rect 42166 30742 42230 30806
rect 34278 30606 34342 30670
rect 34006 30470 34070 30534
rect 42846 30470 42910 30534
rect 37406 29926 37470 29990
rect 34142 29110 34206 29174
rect 34278 28974 34342 29038
rect 1230 28838 1294 28902
rect 42166 28838 42230 28902
rect 34006 27750 34070 27814
rect 34414 27614 34478 27678
rect 1230 27342 1294 27406
rect 42166 27342 42230 27406
rect 8846 26662 8910 26726
rect 34278 26390 34342 26454
rect 8574 26254 8638 26318
rect 34142 26254 34206 26318
rect 20134 25710 20198 25774
rect 20950 25710 21014 25774
rect 21494 25710 21558 25774
rect 22174 25710 22238 25774
rect 22718 25710 22782 25774
rect 23398 25710 23462 25774
rect 1230 25574 1294 25638
rect 8982 25302 9046 25366
rect 19318 25438 19382 25502
rect 20134 25438 20198 25502
rect 20406 25438 20470 25502
rect 20678 25438 20742 25502
rect 20950 25438 21014 25502
rect 21494 25438 21558 25502
rect 21630 25438 21694 25502
rect 21902 25438 21966 25502
rect 22174 25438 22238 25502
rect 22718 25438 22782 25502
rect 22854 25438 22918 25502
rect 23126 25438 23190 25502
rect 23398 25438 23462 25502
rect 23942 25166 24006 25230
rect 24214 25438 24278 25502
rect 42166 25438 42230 25502
rect 21494 24894 21558 24958
rect 22582 24894 22646 24958
rect 34414 24894 34478 24958
rect 34278 24758 34342 24822
rect 41622 24758 41686 24822
rect 8846 24078 8910 24142
rect 1230 23806 1294 23870
rect 19590 24078 19654 24142
rect 21494 24214 21558 24278
rect 22582 24214 22646 24278
rect 8846 23806 8910 23870
rect 41622 23942 41686 24006
rect 42166 23806 42230 23870
rect 34142 23534 34206 23598
rect 19726 23398 19790 23462
rect 23942 23398 24006 23462
rect 40126 23398 40190 23462
rect 42846 23398 42910 23462
rect 40793 23034 40857 23098
rect 8982 22582 9046 22646
rect 12246 22446 12310 22510
rect 1230 22174 1294 22238
rect 19590 22310 19654 22374
rect 19590 22174 19654 22238
rect 20270 22174 20334 22238
rect 20814 22174 20878 22238
rect 22038 22174 22102 22238
rect 22718 22174 22782 22238
rect 23262 22174 23326 22238
rect 24078 22174 24142 22238
rect 24350 22174 24414 22238
rect 34278 22174 34342 22238
rect 42166 22174 42230 22238
rect 19590 21766 19654 21830
rect 20270 21766 20334 21830
rect 18094 21630 18158 21694
rect 20814 21766 20878 21830
rect 22038 21766 22102 21830
rect 22718 21766 22782 21830
rect 23262 21766 23326 21830
rect 24078 21766 24142 21830
rect 24350 21766 24414 21830
rect 26254 21630 26318 21694
rect 19726 21494 19790 21558
rect 26254 21358 26318 21422
rect 8846 21222 8910 21286
rect 10478 21086 10542 21150
rect 27886 21222 27950 21286
rect 28022 21222 28086 21286
rect 3950 20814 4014 20878
rect 14150 20678 14214 20742
rect 14694 20678 14758 20742
rect 14966 20678 15030 20742
rect 18094 20814 18158 20878
rect 15238 20678 15302 20742
rect 27886 20814 27950 20878
rect 28022 20814 28086 20878
rect 28022 20678 28086 20742
rect 28702 20678 28766 20742
rect 28974 20678 29038 20742
rect 29382 20678 29446 20742
rect 40126 20678 40190 20742
rect 1230 20406 1294 20470
rect 14150 20406 14214 20470
rect 2641 20341 2705 20345
rect 2641 20285 2645 20341
rect 2645 20285 2701 20341
rect 2701 20285 2705 20341
rect 2641 20281 2705 20285
rect 14150 20270 14214 20334
rect 14694 20406 14758 20470
rect 14694 20270 14758 20334
rect 14966 20406 15030 20470
rect 14966 20270 15030 20334
rect 15238 20406 15302 20470
rect 15238 20270 15302 20334
rect 28022 20406 28086 20470
rect 28022 20270 28086 20334
rect 28702 20406 28766 20470
rect 28702 20270 28766 20334
rect 28974 20406 29038 20470
rect 28974 20270 29038 20334
rect 29382 20406 29446 20470
rect 42166 20406 42230 20470
rect 29246 20270 29310 20334
rect 14150 19998 14214 20062
rect 14150 19862 14214 19926
rect 14694 19998 14758 20062
rect 14558 19862 14622 19926
rect 14966 19998 15030 20062
rect 15102 19862 15166 19926
rect 15238 19998 15302 20062
rect 15238 19862 15302 19926
rect 28022 19998 28086 20062
rect 2454 19454 2518 19518
rect 14150 19590 14214 19654
rect 14150 19454 14214 19518
rect 14558 19590 14622 19654
rect 14558 19454 14622 19518
rect 15102 19590 15166 19654
rect 14966 19454 15030 19518
rect 15238 19590 15302 19654
rect 15238 19454 15302 19518
rect 28294 19862 28358 19926
rect 28702 19998 28766 20062
rect 28430 19862 28494 19926
rect 28974 19998 29038 20062
rect 28838 19862 28902 19926
rect 29246 19998 29310 20062
rect 29246 19862 29310 19926
rect 28294 19590 28358 19654
rect 28158 19454 28222 19518
rect 28430 19590 28494 19654
rect 28430 19454 28494 19518
rect 28838 19590 28902 19654
rect 28838 19454 28902 19518
rect 29246 19590 29310 19654
rect 29246 19454 29310 19518
rect 14150 19182 14214 19246
rect 14558 19182 14622 19246
rect 14966 19182 15030 19246
rect 14966 19046 15030 19110
rect 15238 19182 15302 19246
rect 15238 19046 15302 19110
rect 1230 18910 1294 18974
rect 2454 18910 2518 18974
rect 28158 19182 28222 19246
rect 28022 19046 28086 19110
rect 28430 19182 28494 19246
rect 28430 19046 28494 19110
rect 28838 19182 28902 19246
rect 25166 18910 25230 18974
rect 14966 18774 15030 18838
rect 15102 18638 15166 18702
rect 15238 18774 15302 18838
rect 15374 18638 15438 18702
rect 12246 18502 12310 18566
rect 3950 18230 4014 18294
rect 11838 18230 11902 18294
rect 12246 18230 12310 18294
rect 12382 18230 12446 18294
rect 12518 18230 12582 18294
rect 15782 18502 15846 18566
rect 15102 18366 15166 18430
rect 15374 18366 15438 18430
rect 18230 18366 18294 18430
rect 16190 18230 16254 18294
rect 550 18094 614 18158
rect 3814 18094 3878 18158
rect 14150 17958 14214 18022
rect 14694 17958 14758 18022
rect 15782 17958 15846 18022
rect 16190 17958 16254 18022
rect 18230 18094 18294 18158
rect 10478 17686 10542 17750
rect 11838 17686 11902 17750
rect 12382 17686 12446 17750
rect 12518 17686 12582 17750
rect 12246 17414 12310 17478
rect 12654 17414 12718 17478
rect 14150 17686 14214 17750
rect 14150 17550 14214 17614
rect 14694 17686 14758 17750
rect 14694 17550 14758 17614
rect 13062 17414 13126 17478
rect 1230 17142 1294 17206
rect 14150 17278 14214 17342
rect 14694 17278 14758 17342
rect 3270 17142 3334 17206
rect 14286 17142 14350 17206
rect 14694 17142 14758 17206
rect 15102 17142 15166 17206
rect 18366 17686 18430 17750
rect 25166 18638 25230 18702
rect 28022 18774 28086 18838
rect 28158 18638 28222 18702
rect 28430 18774 28494 18838
rect 28702 18638 28766 18702
rect 27886 18502 27950 18566
rect 28158 18366 28222 18430
rect 27614 18230 27678 18294
rect 28702 18366 28766 18430
rect 29246 19182 29310 19246
rect 41622 19182 41686 19246
rect 41622 18910 41686 18974
rect 42166 18910 42230 18974
rect 30470 18230 30534 18294
rect 31150 18230 31214 18294
rect 31694 18230 31758 18294
rect 26526 17958 26590 18022
rect 27614 17958 27678 18022
rect 27886 17958 27950 18022
rect 28974 17958 29038 18022
rect 29246 17958 29310 18022
rect 42846 17822 42910 17886
rect 25302 17686 25366 17750
rect 26526 17686 26590 17750
rect 18366 17414 18430 17478
rect 15238 17142 15302 17206
rect 18366 17278 18430 17342
rect 25302 17414 25366 17478
rect 28974 17686 29038 17750
rect 28974 17550 29038 17614
rect 29246 17686 29310 17750
rect 29246 17550 29310 17614
rect 30470 17686 30534 17750
rect 30470 17414 30534 17478
rect 31150 17686 31214 17750
rect 31694 17686 31758 17750
rect 30878 17414 30942 17478
rect 39854 17686 39918 17750
rect 25302 17278 25366 17342
rect 28158 17142 28222 17206
rect 28702 17142 28766 17206
rect 28974 17278 29038 17342
rect 28974 17142 29038 17206
rect 29246 17278 29310 17342
rect 29246 17142 29310 17206
rect 41622 17142 41686 17206
rect 42166 17142 42230 17206
rect 18366 17006 18430 17070
rect 14286 16870 14350 16934
rect 3270 16734 3334 16798
rect 14150 16734 14214 16798
rect 14694 16870 14758 16934
rect 14558 16734 14622 16798
rect 15102 16870 15166 16934
rect 15102 16734 15166 16798
rect 15238 16870 15302 16934
rect 25302 17006 25366 17070
rect 15510 16734 15574 16798
rect 14150 16462 14214 16526
rect 14286 16326 14350 16390
rect 14558 16462 14622 16526
rect 14694 16326 14758 16390
rect 15102 16462 15166 16526
rect 15102 16326 15166 16390
rect 15510 16462 15574 16526
rect 15510 16326 15574 16390
rect 28158 16870 28222 16934
rect 28158 16734 28222 16798
rect 28702 16870 28766 16934
rect 28566 16734 28630 16798
rect 28974 16870 29038 16934
rect 28974 16734 29038 16798
rect 29246 16870 29310 16934
rect 29246 16734 29310 16798
rect 28158 16462 28222 16526
rect 28294 16326 28358 16390
rect 28566 16462 28630 16526
rect 28566 16326 28630 16390
rect 28974 16462 29038 16526
rect 28974 16326 29038 16390
rect 29246 16462 29310 16526
rect 29246 16326 29310 16390
rect 41622 16462 41686 16526
rect 11974 15918 12038 15982
rect 12246 15918 12310 15982
rect 12654 16054 12718 16118
rect 12790 15918 12854 15982
rect 13062 16054 13126 16118
rect 14286 16054 14350 16118
rect 14286 15918 14350 15982
rect 14694 16054 14758 16118
rect 15102 16054 15166 16118
rect 14694 15918 14758 15982
rect 14966 15918 15030 15982
rect 15510 16054 15574 16118
rect 15510 15918 15574 15982
rect 28294 16054 28358 16118
rect 28158 15918 28222 15982
rect 28566 16054 28630 16118
rect 28566 15918 28630 15982
rect 28974 16054 29038 16118
rect 29246 16054 29310 16118
rect 30470 16054 30534 16118
rect 28974 15918 29038 15982
rect 29382 15918 29446 15982
rect 30878 16054 30942 16118
rect 31014 15918 31078 15982
rect 31286 15918 31350 15982
rect 12790 15646 12854 15710
rect 14286 15646 14350 15710
rect 1230 15510 1294 15574
rect 14150 15510 14214 15574
rect 14694 15646 14758 15710
rect 14694 15510 14758 15574
rect 14966 15646 15030 15710
rect 14966 15510 15030 15574
rect 15510 15646 15574 15710
rect 15238 15510 15302 15574
rect 28158 15646 28222 15710
rect 28022 15510 28086 15574
rect 28566 15646 28630 15710
rect 28566 15510 28630 15574
rect 28974 15646 29038 15710
rect 28974 15510 29038 15574
rect 29382 15646 29446 15710
rect 29246 15510 29310 15574
rect 3814 15374 3878 15438
rect 3406 15238 3470 15302
rect 11974 15238 12038 15302
rect 10478 15102 10542 15166
rect 10886 15102 10950 15166
rect 12246 15238 12310 15302
rect 12110 15102 12174 15166
rect 12518 15102 12582 15166
rect 14150 15238 14214 15302
rect 14694 15238 14758 15302
rect 14966 15238 15030 15302
rect 15238 15238 15302 15302
rect 15374 15102 15438 15166
rect 18230 14966 18294 15030
rect 12110 14830 12174 14894
rect 12518 14830 12582 14894
rect 42166 15374 42230 15438
rect 28022 15238 28086 15302
rect 28566 15238 28630 15302
rect 28974 15238 29038 15302
rect 29246 15238 29310 15302
rect 31014 15238 31078 15302
rect 31286 15238 31350 15302
rect 32782 15102 32846 15166
rect 34686 15102 34750 15166
rect 39854 15102 39918 15166
rect 34686 14830 34750 14894
rect 15374 14694 15438 14758
rect 19590 14694 19654 14758
rect 25166 14694 25230 14758
rect 40126 14830 40190 14894
rect 34686 14694 34750 14758
rect 17686 14558 17750 14622
rect 18230 14558 18294 14622
rect 17686 14286 17750 14350
rect 19046 14150 19110 14214
rect 20814 14150 20878 14214
rect 21494 14150 21558 14214
rect 22038 14150 22102 14214
rect 22718 14150 22782 14214
rect 23126 14150 23190 14214
rect 23262 14150 23326 14214
rect 23806 14150 23870 14214
rect 23942 14150 24006 14214
rect 1230 13742 1294 13806
rect 10478 14014 10542 14078
rect 9526 13742 9590 13806
rect 19046 13742 19110 13806
rect 20814 13742 20878 13806
rect 21494 13742 21558 13806
rect 22038 13742 22102 13806
rect 22718 13742 22782 13806
rect 22582 13606 22646 13670
rect 23126 13742 23190 13806
rect 23262 13742 23326 13806
rect 23806 13742 23870 13806
rect 23942 13742 24006 13806
rect 42166 13742 42230 13806
rect 32782 13470 32846 13534
rect 34822 13334 34886 13398
rect 2641 12874 2705 12938
rect 40793 12859 40857 12863
rect 40793 12803 40797 12859
rect 40797 12803 40853 12859
rect 40853 12803 40857 12859
rect 40793 12799 40857 12803
rect 3406 12518 3470 12582
rect 4086 12382 4150 12446
rect 10886 12518 10950 12582
rect 19590 12518 19654 12582
rect 20134 12518 20198 12582
rect 25166 12518 25230 12582
rect 9390 12382 9454 12446
rect 1230 12246 1294 12310
rect 40126 12246 40190 12310
rect 34686 12110 34750 12174
rect 20270 11702 20334 11766
rect 22582 11838 22646 11902
rect 42166 12246 42230 12310
rect 34686 11838 34750 11902
rect 3270 11022 3334 11086
rect 9526 11158 9590 11222
rect 9526 11022 9590 11086
rect 20270 11022 20334 11086
rect 19998 10886 20062 10950
rect 19726 10750 19790 10814
rect 20950 10750 21014 10814
rect 3270 10478 3334 10542
rect 20134 10614 20198 10678
rect 22446 10750 22510 10814
rect 20134 10478 20198 10542
rect 20270 10478 20334 10542
rect 21494 10478 21558 10542
rect 21630 10478 21694 10542
rect 22174 10478 22238 10542
rect 22718 10478 22782 10542
rect 22854 10478 22918 10542
rect 23670 10750 23734 10814
rect 23398 10478 23462 10542
rect 23942 10478 24006 10542
rect 24078 10478 24142 10542
rect 34822 10614 34886 10678
rect 1230 10342 1294 10406
rect 42166 10342 42230 10406
rect 23398 10206 23462 10270
rect 21494 10070 21558 10134
rect 20134 9934 20198 9998
rect 4086 9662 4150 9726
rect 9390 9662 9454 9726
rect 20134 9662 20198 9726
rect 20814 9662 20878 9726
rect 22174 9934 22238 9998
rect 22718 9934 22782 9998
rect 23942 9934 24006 9998
rect 23262 9662 23326 9726
rect 9390 9526 9454 9590
rect 19998 9526 20062 9590
rect 20678 9254 20742 9318
rect 34686 9254 34750 9318
rect 20134 9118 20198 9182
rect 20814 9118 20878 9182
rect 23262 9118 23326 9182
rect 1230 8846 1294 8910
rect 3270 8710 3334 8774
rect 19046 8710 19110 8774
rect 24486 8710 24550 8774
rect 42166 8710 42230 8774
rect 19318 8438 19382 8502
rect 20678 8438 20742 8502
rect 24350 8438 24414 8502
rect 3270 8302 3334 8366
rect 9526 8302 9590 8366
rect 9526 8166 9590 8230
rect 19318 8030 19382 8094
rect 24350 8030 24414 8094
rect 1230 7078 1294 7142
rect 42166 7078 42230 7142
rect 9390 6942 9454 7006
rect 19046 6942 19110 7006
rect 24486 6942 24550 7006
rect 9526 6670 9590 6734
rect 550 5582 614 5646
rect 1230 5310 1294 5374
rect 9390 5446 9454 5510
rect 9254 5310 9318 5374
rect 42166 5310 42230 5374
rect 9526 4086 9590 4150
rect 9390 3950 9454 4014
rect 1230 3814 1294 3878
rect 42166 3814 42230 3878
rect 5990 3134 6054 3198
rect 10750 3134 10814 3198
rect 12110 3134 12174 3198
rect 13198 3192 13262 3198
rect 13198 3136 13228 3192
rect 13228 3136 13262 3192
rect 13198 3134 13262 3136
rect 14422 3134 14486 3198
rect 15510 3192 15574 3198
rect 15510 3136 15564 3192
rect 15564 3136 15574 3192
rect 15510 3134 15574 3136
rect 16734 3134 16798 3198
rect 17958 3134 18022 3198
rect 19046 3192 19110 3198
rect 19046 3136 19068 3192
rect 19068 3136 19110 3192
rect 19046 3134 19110 3136
rect 20270 3134 20334 3198
rect 21358 3192 21422 3198
rect 21358 3136 21404 3192
rect 21404 3136 21422 3192
rect 21358 3134 21422 3136
rect 22582 3134 22646 3198
rect 23806 3134 23870 3198
rect 9254 2590 9318 2654
rect 550 2454 614 2518
rect 9526 2454 9590 2518
rect 2046 2046 2110 2110
rect 42166 2046 42230 2110
rect 2046 1788 2110 1838
rect 2046 1774 2066 1788
rect 2066 1774 2110 1788
rect 2182 1638 2246 1702
rect 3814 1638 3878 1702
rect 5446 1638 5510 1702
rect 7078 1638 7142 1702
rect 9390 1774 9454 1838
rect 8710 1638 8774 1702
rect 10342 1638 10406 1702
rect 12246 1638 12310 1702
rect 13742 1638 13806 1702
rect 15374 1638 15438 1702
rect 17278 1638 17342 1702
rect 18774 1638 18838 1702
rect 20678 1638 20742 1702
rect 22310 1638 22374 1702
rect 23534 1638 23598 1702
rect 25438 1638 25502 1702
rect 27342 1638 27406 1702
rect 28974 1638 29038 1702
rect 30606 1638 30670 1702
rect 32238 1638 32302 1702
rect 34006 1638 34070 1702
rect 35638 1638 35702 1702
rect 37406 1638 37470 1702
rect 39038 1638 39102 1702
rect 40806 1638 40870 1702
rect 958 1230 1022 1294
rect 1094 1230 1158 1294
rect 1230 1230 1294 1294
rect 2182 1230 2246 1294
rect 3814 1230 3878 1294
rect 5446 1230 5510 1294
rect 7078 1230 7142 1294
rect 8710 1230 8774 1294
rect 10342 1230 10406 1294
rect 12246 1230 12310 1294
rect 13742 1230 13806 1294
rect 15374 1230 15438 1294
rect 17278 1230 17342 1294
rect 18774 1230 18838 1294
rect 20678 1230 20742 1294
rect 22310 1230 22374 1294
rect 23534 1230 23598 1294
rect 25438 1230 25502 1294
rect 27342 1230 27406 1294
rect 28974 1230 29038 1294
rect 30606 1230 30670 1294
rect 32238 1230 32302 1294
rect 34006 1230 34070 1294
rect 35638 1230 35702 1294
rect 37406 1230 37470 1294
rect 39038 1230 39102 1294
rect 40806 1230 40870 1294
rect 42166 1230 42230 1294
rect 42302 1230 42366 1294
rect 42438 1230 42502 1294
rect 958 1094 1022 1158
rect 1094 1094 1158 1158
rect 1230 1094 1294 1158
rect 42166 1094 42230 1158
rect 42302 1094 42366 1158
rect 42438 1094 42502 1158
rect 958 958 1022 1022
rect 1094 958 1158 1022
rect 1230 958 1294 1022
rect 42166 958 42230 1022
rect 42302 958 42366 1022
rect 42438 958 42502 1022
rect 278 550 342 614
rect 414 550 478 614
rect 550 550 614 614
rect 9526 550 9590 614
rect 42846 550 42910 614
rect 42982 550 43046 614
rect 43118 550 43182 614
rect 278 414 342 478
rect 414 414 478 478
rect 550 414 614 478
rect 42846 414 42910 478
rect 42982 414 43046 478
rect 43118 414 43182 478
rect 278 278 342 342
rect 414 278 478 342
rect 550 278 614 342
rect 42846 278 42910 342
rect 42982 278 43046 342
rect 43118 278 43182 342
<< metal4 >>
rect 272 32846 620 32852
rect 272 32782 278 32846
rect 342 32782 414 32846
rect 478 32782 550 32846
rect 614 32782 620 32846
rect 272 32710 620 32782
rect 272 32646 278 32710
rect 342 32646 414 32710
rect 478 32646 550 32710
rect 614 32646 620 32710
rect 272 32574 620 32646
rect 272 32510 278 32574
rect 342 32510 414 32574
rect 478 32510 550 32574
rect 614 32510 620 32574
rect 272 18158 620 32510
rect 272 18094 550 18158
rect 614 18094 620 18158
rect 272 5646 620 18094
rect 272 5582 550 5646
rect 614 5582 620 5646
rect 272 2518 620 5582
rect 272 2454 550 2518
rect 614 2454 620 2518
rect 272 614 620 2454
rect 952 32166 1300 32172
rect 952 32102 958 32166
rect 1022 32102 1094 32166
rect 1158 32102 1230 32166
rect 1294 32102 1300 32166
rect 952 32030 1300 32102
rect 952 31966 958 32030
rect 1022 31966 1094 32030
rect 1158 31966 1230 32030
rect 1294 31966 1300 32030
rect 952 31894 1300 31966
rect 952 31830 958 31894
rect 1022 31830 1094 31894
rect 1158 31830 1230 31894
rect 1294 31830 1300 31894
rect 952 30806 1300 31830
rect 2176 31894 2252 31900
rect 2176 31830 2182 31894
rect 2246 31830 2252 31894
rect 2176 31486 2252 31830
rect 2176 31454 2182 31486
rect 2181 31422 2182 31454
rect 2246 31454 2252 31486
rect 3808 31894 3884 31900
rect 3808 31830 3814 31894
rect 3878 31830 3884 31894
rect 3808 31486 3884 31830
rect 3808 31454 3814 31486
rect 2246 31422 2247 31454
rect 2181 31421 2247 31422
rect 3813 31422 3814 31454
rect 3878 31454 3884 31486
rect 5304 31894 5380 31900
rect 5304 31830 5310 31894
rect 5374 31830 5380 31894
rect 5304 31486 5380 31830
rect 5304 31454 5310 31486
rect 3878 31422 3879 31454
rect 3813 31421 3879 31422
rect 5309 31422 5310 31454
rect 5374 31454 5380 31486
rect 7072 31894 7148 31900
rect 7072 31830 7078 31894
rect 7142 31830 7148 31894
rect 7072 31486 7148 31830
rect 7072 31454 7078 31486
rect 5374 31422 5375 31454
rect 5309 31421 5375 31422
rect 7077 31422 7078 31454
rect 7142 31454 7148 31486
rect 7142 31422 7143 31454
rect 7077 31421 7143 31422
rect 952 30742 1230 30806
rect 1294 30742 1300 30806
rect 952 28902 1300 30742
rect 952 28838 1230 28902
rect 1294 28838 1300 28902
rect 952 27406 1300 28838
rect 952 27342 1230 27406
rect 1294 27342 1300 27406
rect 952 25638 1300 27342
rect 8568 26318 8644 33124
rect 8704 31894 8780 31900
rect 8704 31830 8710 31894
rect 8774 31830 8780 31894
rect 8704 31486 8780 31830
rect 8704 31454 8710 31486
rect 8709 31422 8710 31454
rect 8774 31454 8780 31486
rect 10336 31894 10412 31900
rect 10336 31830 10342 31894
rect 10406 31830 10412 31894
rect 10336 31486 10412 31830
rect 10336 31454 10342 31486
rect 8774 31422 8775 31454
rect 8709 31421 8775 31422
rect 10341 31422 10342 31454
rect 10406 31454 10412 31486
rect 12104 31894 12180 31900
rect 12104 31830 12110 31894
rect 12174 31830 12180 31894
rect 12104 31486 12180 31830
rect 12104 31454 12110 31486
rect 10406 31422 10407 31454
rect 10341 31421 10407 31422
rect 12109 31422 12110 31454
rect 12174 31454 12180 31486
rect 13736 31894 13812 31900
rect 13736 31830 13742 31894
rect 13806 31830 13812 31894
rect 13736 31486 13812 31830
rect 13736 31454 13742 31486
rect 12174 31422 12175 31454
rect 12109 31421 12175 31422
rect 13741 31422 13742 31454
rect 13806 31454 13812 31486
rect 15640 31894 15716 31900
rect 15640 31830 15646 31894
rect 15710 31830 15716 31894
rect 15640 31486 15716 31830
rect 15640 31454 15646 31486
rect 13806 31422 13807 31454
rect 13741 31421 13807 31422
rect 15645 31422 15646 31454
rect 15710 31454 15716 31486
rect 17272 31894 17348 31900
rect 17272 31830 17278 31894
rect 17342 31830 17348 31894
rect 17272 31486 17348 31830
rect 17272 31454 17278 31486
rect 15710 31422 15711 31454
rect 15645 31421 15711 31422
rect 17277 31422 17278 31454
rect 17342 31454 17348 31486
rect 18768 31894 18844 31900
rect 18768 31830 18774 31894
rect 18838 31830 18844 31894
rect 18768 31486 18844 31830
rect 18768 31454 18774 31486
rect 17342 31422 17343 31454
rect 17277 31421 17343 31422
rect 18773 31422 18774 31454
rect 18838 31454 18844 31486
rect 18838 31422 18839 31454
rect 18773 31421 18839 31422
rect 8568 26286 8574 26318
rect 8573 26254 8574 26286
rect 8638 26286 8644 26318
rect 8840 26726 8916 26732
rect 8840 26662 8846 26726
rect 8910 26662 8916 26726
rect 8638 26254 8639 26286
rect 8573 26253 8639 26254
rect 952 25574 1230 25638
rect 1294 25574 1300 25638
rect 952 23870 1300 25574
rect 8840 24142 8916 26662
rect 19312 25502 19388 33124
rect 20264 31894 20340 31900
rect 20264 31830 20270 31894
rect 20334 31830 20340 31894
rect 20264 31486 20340 31830
rect 20264 31454 20270 31486
rect 20269 31422 20270 31454
rect 20334 31454 20340 31486
rect 20334 31422 20335 31454
rect 20269 31421 20335 31422
rect 19312 25470 19318 25502
rect 19317 25438 19318 25470
rect 19382 25470 19388 25502
rect 20128 25774 20204 25780
rect 20128 25710 20134 25774
rect 20198 25710 20204 25774
rect 20128 25502 20204 25710
rect 20128 25470 20134 25502
rect 19382 25438 19383 25470
rect 19317 25437 19383 25438
rect 20133 25438 20134 25470
rect 20198 25470 20204 25502
rect 20400 25502 20476 33124
rect 20400 25470 20406 25502
rect 20198 25438 20199 25470
rect 20133 25437 20199 25438
rect 20405 25438 20406 25470
rect 20470 25470 20476 25502
rect 20672 25502 20748 33124
rect 20949 25774 21015 25775
rect 20949 25742 20950 25774
rect 20672 25470 20678 25502
rect 20470 25438 20471 25470
rect 20405 25437 20471 25438
rect 20677 25438 20678 25470
rect 20742 25470 20748 25502
rect 20944 25710 20950 25742
rect 21014 25742 21015 25774
rect 21488 25774 21564 25780
rect 21014 25710 21020 25742
rect 20944 25502 21020 25710
rect 20742 25438 20743 25470
rect 20677 25437 20743 25438
rect 20944 25438 20950 25502
rect 21014 25438 21020 25502
rect 21488 25710 21494 25774
rect 21558 25710 21564 25774
rect 21488 25502 21564 25710
rect 21488 25470 21494 25502
rect 20944 25432 21020 25438
rect 21493 25438 21494 25470
rect 21558 25470 21564 25502
rect 21624 25502 21700 33124
rect 21624 25470 21630 25502
rect 21558 25438 21559 25470
rect 21493 25437 21559 25438
rect 21629 25438 21630 25470
rect 21694 25470 21700 25502
rect 21896 25502 21972 33124
rect 22304 31894 22380 31900
rect 22304 31830 22310 31894
rect 22374 31830 22380 31894
rect 22304 31486 22380 31830
rect 22304 31454 22310 31486
rect 22309 31422 22310 31454
rect 22374 31454 22380 31486
rect 22374 31422 22375 31454
rect 22309 31421 22375 31422
rect 22173 25774 22239 25775
rect 22173 25742 22174 25774
rect 21896 25470 21902 25502
rect 21694 25438 21695 25470
rect 21629 25437 21695 25438
rect 21901 25438 21902 25470
rect 21966 25470 21972 25502
rect 22168 25710 22174 25742
rect 22238 25742 22239 25774
rect 22712 25774 22788 25780
rect 22238 25710 22244 25742
rect 22168 25502 22244 25710
rect 21966 25438 21967 25470
rect 21901 25437 21967 25438
rect 22168 25438 22174 25502
rect 22238 25438 22244 25502
rect 22712 25710 22718 25774
rect 22782 25710 22788 25774
rect 22712 25502 22788 25710
rect 22712 25470 22718 25502
rect 22168 25432 22244 25438
rect 22717 25438 22718 25470
rect 22782 25470 22788 25502
rect 22848 25502 22924 33124
rect 22848 25470 22854 25502
rect 22782 25438 22783 25470
rect 22717 25437 22783 25438
rect 22853 25438 22854 25470
rect 22918 25470 22924 25502
rect 23120 25502 23196 33124
rect 23800 31894 23876 31900
rect 23800 31830 23806 31894
rect 23870 31830 23876 31894
rect 23800 31486 23876 31830
rect 23800 31454 23806 31486
rect 23805 31422 23806 31454
rect 23870 31454 23876 31486
rect 23870 31422 23871 31454
rect 23805 31421 23871 31422
rect 23397 25774 23463 25775
rect 23397 25742 23398 25774
rect 23120 25470 23126 25502
rect 22918 25438 22919 25470
rect 22853 25437 22919 25438
rect 23125 25438 23126 25470
rect 23190 25470 23196 25502
rect 23392 25710 23398 25742
rect 23462 25742 23463 25774
rect 23462 25710 23468 25742
rect 23392 25502 23468 25710
rect 23190 25438 23191 25470
rect 23125 25437 23191 25438
rect 23392 25438 23398 25502
rect 23462 25438 23468 25502
rect 24208 25502 24284 33124
rect 34272 32574 34348 32580
rect 34272 32510 34278 32574
rect 34342 32510 34348 32574
rect 25568 31894 25644 31900
rect 25568 31830 25574 31894
rect 25638 31830 25644 31894
rect 25568 31486 25644 31830
rect 25568 31454 25574 31486
rect 25573 31422 25574 31454
rect 25638 31454 25644 31486
rect 27200 31894 27276 31900
rect 27200 31830 27206 31894
rect 27270 31830 27276 31894
rect 27200 31486 27276 31830
rect 27200 31454 27206 31486
rect 25638 31422 25639 31454
rect 25573 31421 25639 31422
rect 27205 31422 27206 31454
rect 27270 31454 27276 31486
rect 28968 31894 29044 31900
rect 28968 31830 28974 31894
rect 29038 31830 29044 31894
rect 28968 31486 29044 31830
rect 28968 31454 28974 31486
rect 27270 31422 27271 31454
rect 27205 31421 27271 31422
rect 28973 31422 28974 31454
rect 29038 31454 29044 31486
rect 30600 31894 30676 31900
rect 30600 31830 30606 31894
rect 30670 31830 30676 31894
rect 30600 31486 30676 31830
rect 30600 31454 30606 31486
rect 29038 31422 29039 31454
rect 28973 31421 29039 31422
rect 30605 31422 30606 31454
rect 30670 31454 30676 31486
rect 32232 31894 32308 31900
rect 32232 31830 32238 31894
rect 32302 31830 32308 31894
rect 32232 31486 32308 31830
rect 32232 31454 32238 31486
rect 30670 31422 30671 31454
rect 30605 31421 30671 31422
rect 32237 31422 32238 31454
rect 32302 31454 32308 31486
rect 34000 31894 34076 31900
rect 34000 31830 34006 31894
rect 34070 31830 34076 31894
rect 34000 31486 34076 31830
rect 34000 31454 34006 31486
rect 32302 31422 32303 31454
rect 32237 31421 32303 31422
rect 34005 31422 34006 31454
rect 34070 31454 34076 31486
rect 34070 31422 34071 31454
rect 34005 31421 34071 31422
rect 34141 31350 34207 31351
rect 34141 31318 34142 31350
rect 34136 31286 34142 31318
rect 34206 31318 34207 31350
rect 34206 31286 34212 31318
rect 34005 30534 34071 30535
rect 34005 30502 34006 30534
rect 34000 30470 34006 30502
rect 34070 30502 34071 30534
rect 34070 30470 34076 30502
rect 34000 27814 34076 30470
rect 34136 29174 34212 31286
rect 34272 30670 34348 32510
rect 35632 31894 35708 31900
rect 35632 31830 35638 31894
rect 35702 31830 35708 31894
rect 35632 31486 35708 31830
rect 35632 31454 35638 31486
rect 35637 31422 35638 31454
rect 35702 31454 35708 31486
rect 37264 31894 37340 31900
rect 37264 31830 37270 31894
rect 37334 31830 37340 31894
rect 37264 31486 37340 31830
rect 37264 31454 37270 31486
rect 35702 31422 35703 31454
rect 35637 31421 35703 31422
rect 37269 31422 37270 31454
rect 37334 31454 37340 31486
rect 37334 31422 37335 31454
rect 37269 31421 37335 31422
rect 34272 30638 34278 30670
rect 34277 30606 34278 30638
rect 34342 30638 34348 30670
rect 34342 30606 34343 30638
rect 34277 30605 34343 30606
rect 37400 29990 37476 33124
rect 42840 32846 43188 32852
rect 42840 32782 42846 32846
rect 42910 32782 42982 32846
rect 43046 32782 43118 32846
rect 43182 32782 43188 32846
rect 42840 32710 43188 32782
rect 42840 32646 42846 32710
rect 42910 32646 42982 32710
rect 43046 32646 43118 32710
rect 43182 32646 43188 32710
rect 42840 32574 43188 32646
rect 42840 32510 42846 32574
rect 42910 32510 42982 32574
rect 43046 32510 43118 32574
rect 43182 32510 43188 32574
rect 42160 32166 42508 32172
rect 42160 32102 42166 32166
rect 42230 32102 42302 32166
rect 42366 32102 42438 32166
rect 42502 32102 42508 32166
rect 42160 32030 42508 32102
rect 42160 31966 42166 32030
rect 42230 31966 42302 32030
rect 42366 31966 42438 32030
rect 42502 31966 42508 32030
rect 38896 31894 38972 31900
rect 38896 31830 38902 31894
rect 38966 31830 38972 31894
rect 38896 31486 38972 31830
rect 38896 31454 38902 31486
rect 38901 31422 38902 31454
rect 38966 31454 38972 31486
rect 40664 31894 40740 31900
rect 40664 31830 40670 31894
rect 40734 31830 40740 31894
rect 40664 31486 40740 31830
rect 40664 31454 40670 31486
rect 38966 31422 38967 31454
rect 38901 31421 38967 31422
rect 40669 31422 40670 31454
rect 40734 31454 40740 31486
rect 42160 31894 42508 31966
rect 42160 31830 42166 31894
rect 42230 31830 42302 31894
rect 42366 31830 42438 31894
rect 42502 31830 42508 31894
rect 40734 31422 40735 31454
rect 40669 31421 40735 31422
rect 37400 29958 37406 29990
rect 37405 29926 37406 29958
rect 37470 29958 37476 29990
rect 42160 30806 42508 31830
rect 42160 30742 42166 30806
rect 42230 30742 42508 30806
rect 37470 29926 37471 29958
rect 37405 29925 37471 29926
rect 34136 29110 34142 29174
rect 34206 29110 34212 29174
rect 34136 29104 34212 29110
rect 34000 27750 34006 27814
rect 34070 27750 34076 27814
rect 34000 27744 34076 27750
rect 34272 29038 34348 29044
rect 34272 28974 34278 29038
rect 34342 28974 34348 29038
rect 34272 26454 34348 28974
rect 42160 28902 42508 30742
rect 42160 28838 42166 28902
rect 42230 28838 42508 28902
rect 34272 26422 34278 26454
rect 34277 26390 34278 26422
rect 34342 26422 34348 26454
rect 34408 27678 34484 27684
rect 34408 27614 34414 27678
rect 34478 27614 34484 27678
rect 34342 26390 34343 26422
rect 34277 26389 34343 26390
rect 24208 25470 24214 25502
rect 23392 25432 23468 25438
rect 24213 25438 24214 25470
rect 24278 25470 24284 25502
rect 34136 26318 34212 26324
rect 34136 26254 34142 26318
rect 34206 26254 34212 26318
rect 24278 25438 24279 25470
rect 24213 25437 24279 25438
rect 8840 24110 8846 24142
rect 8845 24078 8846 24110
rect 8910 24110 8916 24142
rect 8976 25366 9052 25372
rect 8976 25302 8982 25366
rect 9046 25302 9052 25366
rect 8910 24078 8911 24110
rect 8845 24077 8911 24078
rect 952 23806 1230 23870
rect 1294 23806 1300 23870
rect 952 22238 1300 23806
rect 952 22174 1230 22238
rect 1294 22174 1300 22238
rect 952 20470 1300 22174
rect 8840 23870 8916 23876
rect 8840 23806 8846 23870
rect 8910 23806 8916 23870
rect 8840 21286 8916 23806
rect 8976 22646 9052 25302
rect 23936 25230 24012 25236
rect 23936 25166 23942 25230
rect 24006 25166 24012 25230
rect 21493 24958 21559 24959
rect 21493 24926 21494 24958
rect 21488 24894 21494 24926
rect 21558 24926 21559 24958
rect 22581 24958 22647 24959
rect 22581 24926 22582 24958
rect 21558 24894 21564 24926
rect 21488 24278 21564 24894
rect 21488 24214 21494 24278
rect 21558 24214 21564 24278
rect 21488 24208 21564 24214
rect 22576 24894 22582 24926
rect 22646 24926 22647 24958
rect 22646 24894 22652 24926
rect 22576 24278 22652 24894
rect 22576 24214 22582 24278
rect 22646 24214 22652 24278
rect 22576 24208 22652 24214
rect 8976 22614 8982 22646
rect 8981 22582 8982 22614
rect 9046 22614 9052 22646
rect 19584 24142 19660 24148
rect 19584 24078 19590 24142
rect 19654 24078 19660 24142
rect 9046 22582 9047 22614
rect 8981 22581 9047 22582
rect 12245 22510 12311 22511
rect 12245 22478 12246 22510
rect 8840 21254 8846 21286
rect 8845 21222 8846 21254
rect 8910 21254 8916 21286
rect 12240 22446 12246 22478
rect 12310 22478 12311 22510
rect 12310 22446 12316 22478
rect 8910 21222 8911 21254
rect 8845 21221 8911 21222
rect 10477 21150 10543 21151
rect 10477 21118 10478 21150
rect 10472 21086 10478 21118
rect 10542 21118 10543 21150
rect 10542 21086 10548 21118
rect 952 20406 1230 20470
rect 1294 20406 1300 20470
rect 952 18974 1300 20406
rect 3944 20878 4020 20884
rect 3944 20814 3950 20878
rect 4014 20814 4020 20878
rect 2640 20345 2706 20346
rect 2640 20281 2641 20345
rect 2705 20281 2706 20345
rect 2640 20280 2706 20281
rect 952 18910 1230 18974
rect 1294 18910 1300 18974
rect 2448 19518 2524 19524
rect 2448 19454 2454 19518
rect 2518 19454 2524 19518
rect 2448 18974 2524 19454
rect 2448 18942 2454 18974
rect 952 17206 1300 18910
rect 2453 18910 2454 18942
rect 2518 18942 2524 18974
rect 2518 18910 2519 18942
rect 2453 18909 2519 18910
rect 952 17142 1230 17206
rect 1294 17142 1300 17206
rect 952 15574 1300 17142
rect 952 15510 1230 15574
rect 1294 15510 1300 15574
rect 952 13806 1300 15510
rect 952 13742 1230 13806
rect 1294 13742 1300 13806
rect 952 12310 1300 13742
rect 2643 12939 2703 20280
rect 3944 18294 4020 20814
rect 3944 18262 3950 18294
rect 3949 18230 3950 18262
rect 4014 18262 4020 18294
rect 4014 18230 4015 18262
rect 3949 18229 4015 18230
rect 3813 18158 3879 18159
rect 3813 18126 3814 18158
rect 3808 18094 3814 18126
rect 3878 18126 3879 18158
rect 3878 18094 3884 18126
rect 3269 17206 3335 17207
rect 3269 17174 3270 17206
rect 3264 17142 3270 17174
rect 3334 17174 3335 17206
rect 3334 17142 3340 17174
rect 3264 16798 3340 17142
rect 3264 16734 3270 16798
rect 3334 16734 3340 16798
rect 3264 16728 3340 16734
rect 3808 15438 3884 18094
rect 10472 17750 10548 21086
rect 12240 18566 12316 22446
rect 19584 22374 19660 24078
rect 19584 22342 19590 22374
rect 19589 22310 19590 22342
rect 19654 22342 19660 22374
rect 19720 23462 19796 23468
rect 19720 23398 19726 23462
rect 19790 23398 19796 23462
rect 23936 23462 24012 25166
rect 34136 23598 34212 26254
rect 34408 24958 34484 27614
rect 34408 24926 34414 24958
rect 34413 24894 34414 24926
rect 34478 24926 34484 24958
rect 42160 27406 42508 28838
rect 42160 27342 42166 27406
rect 42230 27342 42508 27406
rect 42160 25502 42508 27342
rect 42160 25438 42166 25502
rect 42230 25438 42508 25502
rect 34478 24894 34479 24926
rect 34413 24893 34479 24894
rect 34136 23566 34142 23598
rect 34141 23534 34142 23566
rect 34206 23566 34212 23598
rect 34272 24822 34348 24828
rect 34272 24758 34278 24822
rect 34342 24758 34348 24822
rect 41621 24822 41687 24823
rect 41621 24790 41622 24822
rect 34206 23534 34207 23566
rect 34141 23533 34207 23534
rect 23936 23430 23942 23462
rect 19654 22310 19655 22342
rect 19589 22309 19655 22310
rect 19589 22238 19655 22239
rect 19589 22206 19590 22238
rect 19584 22174 19590 22206
rect 19654 22206 19655 22238
rect 19654 22174 19660 22206
rect 19584 21830 19660 22174
rect 19584 21766 19590 21830
rect 19654 21766 19660 21830
rect 19584 21760 19660 21766
rect 18088 21694 18164 21700
rect 18088 21630 18094 21694
rect 18158 21630 18164 21694
rect 18088 20878 18164 21630
rect 19720 21558 19796 23398
rect 23941 23398 23942 23430
rect 24006 23430 24012 23462
rect 24006 23398 24007 23430
rect 23941 23397 24007 23398
rect 20264 22238 20340 22244
rect 20264 22174 20270 22238
rect 20334 22174 20340 22238
rect 20813 22238 20879 22239
rect 20813 22206 20814 22238
rect 20264 21830 20340 22174
rect 20264 21798 20270 21830
rect 20269 21766 20270 21798
rect 20334 21798 20340 21830
rect 20808 22174 20814 22206
rect 20878 22206 20879 22238
rect 22037 22238 22103 22239
rect 22037 22206 22038 22238
rect 20878 22174 20884 22206
rect 20808 21830 20884 22174
rect 20334 21766 20335 21798
rect 20269 21765 20335 21766
rect 20808 21766 20814 21830
rect 20878 21766 20884 21830
rect 20808 21760 20884 21766
rect 22032 22174 22038 22206
rect 22102 22206 22103 22238
rect 22712 22238 22788 22244
rect 22102 22174 22108 22206
rect 22032 21830 22108 22174
rect 22032 21766 22038 21830
rect 22102 21766 22108 21830
rect 22712 22174 22718 22238
rect 22782 22174 22788 22238
rect 23261 22238 23327 22239
rect 23261 22206 23262 22238
rect 22712 21830 22788 22174
rect 22712 21798 22718 21830
rect 22032 21760 22108 21766
rect 22717 21766 22718 21798
rect 22782 21798 22788 21830
rect 23256 22174 23262 22206
rect 23326 22206 23327 22238
rect 24072 22238 24148 22244
rect 23326 22174 23332 22206
rect 23256 21830 23332 22174
rect 22782 21766 22783 21798
rect 22717 21765 22783 21766
rect 23256 21766 23262 21830
rect 23326 21766 23332 21830
rect 24072 22174 24078 22238
rect 24142 22174 24148 22238
rect 24072 21830 24148 22174
rect 24072 21798 24078 21830
rect 23256 21760 23332 21766
rect 24077 21766 24078 21798
rect 24142 21798 24148 21830
rect 24344 22238 24420 22244
rect 24344 22174 24350 22238
rect 24414 22174 24420 22238
rect 34272 22238 34348 24758
rect 41616 24758 41622 24790
rect 41686 24790 41687 24822
rect 41686 24758 41692 24790
rect 41616 24006 41692 24758
rect 41616 23942 41622 24006
rect 41686 23942 41692 24006
rect 41616 23936 41692 23942
rect 42160 23870 42508 25438
rect 42160 23806 42166 23870
rect 42230 23806 42508 23870
rect 40125 23462 40191 23463
rect 40125 23430 40126 23462
rect 34272 22206 34278 22238
rect 24344 21830 24420 22174
rect 34277 22174 34278 22206
rect 34342 22206 34348 22238
rect 40120 23398 40126 23430
rect 40190 23430 40191 23462
rect 40190 23398 40196 23430
rect 34342 22174 34343 22206
rect 34277 22173 34343 22174
rect 24344 21798 24350 21830
rect 24142 21766 24143 21798
rect 24077 21765 24143 21766
rect 24349 21766 24350 21798
rect 24414 21798 24420 21830
rect 24414 21766 24415 21798
rect 24349 21765 24415 21766
rect 26253 21694 26319 21695
rect 26253 21662 26254 21694
rect 19720 21526 19726 21558
rect 19725 21494 19726 21526
rect 19790 21526 19796 21558
rect 26248 21630 26254 21662
rect 26318 21662 26319 21694
rect 26318 21630 26324 21662
rect 19790 21494 19791 21526
rect 19725 21493 19791 21494
rect 26248 21422 26324 21630
rect 26248 21358 26254 21422
rect 26318 21358 26324 21422
rect 26248 21352 26324 21358
rect 27885 21286 27951 21287
rect 27885 21254 27886 21286
rect 18088 20846 18094 20878
rect 18093 20814 18094 20846
rect 18158 20846 18164 20878
rect 27880 21222 27886 21254
rect 27950 21254 27951 21286
rect 28021 21286 28087 21287
rect 28021 21254 28022 21286
rect 27950 21222 27956 21254
rect 27880 20878 27956 21222
rect 18158 20814 18159 20846
rect 18093 20813 18159 20814
rect 27880 20814 27886 20878
rect 27950 20814 27956 20878
rect 27880 20808 27956 20814
rect 28016 21222 28022 21254
rect 28086 21254 28087 21286
rect 28086 21222 28092 21254
rect 28016 20878 28092 21222
rect 28016 20814 28022 20878
rect 28086 20814 28092 20878
rect 28016 20808 28092 20814
rect 14149 20742 14215 20743
rect 14149 20710 14150 20742
rect 14144 20678 14150 20710
rect 14214 20710 14215 20742
rect 14688 20742 14764 20748
rect 14214 20678 14220 20710
rect 14144 20470 14220 20678
rect 14144 20406 14150 20470
rect 14214 20406 14220 20470
rect 14688 20678 14694 20742
rect 14758 20678 14764 20742
rect 14965 20742 15031 20743
rect 14965 20710 14966 20742
rect 14688 20470 14764 20678
rect 14688 20438 14694 20470
rect 14144 20400 14220 20406
rect 14693 20406 14694 20438
rect 14758 20438 14764 20470
rect 14960 20678 14966 20710
rect 15030 20710 15031 20742
rect 15232 20742 15308 20748
rect 15030 20678 15036 20710
rect 14960 20470 15036 20678
rect 14758 20406 14759 20438
rect 14693 20405 14759 20406
rect 14960 20406 14966 20470
rect 15030 20406 15036 20470
rect 15232 20678 15238 20742
rect 15302 20678 15308 20742
rect 28021 20742 28087 20743
rect 28021 20710 28022 20742
rect 15232 20470 15308 20678
rect 15232 20438 15238 20470
rect 14960 20400 15036 20406
rect 15237 20406 15238 20438
rect 15302 20438 15308 20470
rect 28016 20678 28022 20710
rect 28086 20710 28087 20742
rect 28696 20742 28772 20748
rect 28086 20678 28092 20710
rect 28016 20470 28092 20678
rect 15302 20406 15303 20438
rect 15237 20405 15303 20406
rect 28016 20406 28022 20470
rect 28086 20406 28092 20470
rect 28696 20678 28702 20742
rect 28766 20678 28772 20742
rect 28696 20470 28772 20678
rect 28696 20438 28702 20470
rect 28016 20400 28092 20406
rect 28701 20406 28702 20438
rect 28766 20438 28772 20470
rect 28968 20742 29044 20748
rect 28968 20678 28974 20742
rect 29038 20678 29044 20742
rect 28968 20470 29044 20678
rect 28968 20438 28974 20470
rect 28766 20406 28767 20438
rect 28701 20405 28767 20406
rect 28973 20406 28974 20438
rect 29038 20438 29044 20470
rect 29376 20742 29452 20748
rect 29376 20678 29382 20742
rect 29446 20678 29452 20742
rect 29376 20470 29452 20678
rect 40120 20742 40196 23398
rect 40792 23098 40858 23099
rect 40792 23034 40793 23098
rect 40857 23034 40858 23098
rect 40792 23033 40858 23034
rect 40120 20678 40126 20742
rect 40190 20678 40196 20742
rect 40120 20672 40196 20678
rect 29376 20438 29382 20470
rect 29038 20406 29039 20438
rect 28973 20405 29039 20406
rect 29381 20406 29382 20438
rect 29446 20438 29452 20470
rect 29446 20406 29447 20438
rect 29381 20405 29447 20406
rect 14144 20334 14220 20340
rect 14144 20270 14150 20334
rect 14214 20270 14220 20334
rect 14144 20062 14220 20270
rect 14144 20030 14150 20062
rect 14149 19998 14150 20030
rect 14214 20030 14220 20062
rect 14688 20334 14764 20340
rect 14688 20270 14694 20334
rect 14758 20270 14764 20334
rect 14965 20334 15031 20335
rect 14965 20302 14966 20334
rect 14688 20062 14764 20270
rect 14688 20030 14694 20062
rect 14214 19998 14215 20030
rect 14149 19997 14215 19998
rect 14693 19998 14694 20030
rect 14758 20030 14764 20062
rect 14960 20270 14966 20302
rect 15030 20302 15031 20334
rect 15237 20334 15303 20335
rect 15237 20302 15238 20334
rect 15030 20270 15036 20302
rect 14960 20062 15036 20270
rect 14758 19998 14759 20030
rect 14693 19997 14759 19998
rect 14960 19998 14966 20062
rect 15030 19998 15036 20062
rect 14960 19992 15036 19998
rect 15232 20270 15238 20302
rect 15302 20302 15303 20334
rect 28016 20334 28092 20340
rect 15302 20270 15308 20302
rect 15232 20062 15308 20270
rect 15232 19998 15238 20062
rect 15302 19998 15308 20062
rect 28016 20270 28022 20334
rect 28086 20270 28092 20334
rect 28701 20334 28767 20335
rect 28701 20302 28702 20334
rect 28016 20062 28092 20270
rect 28016 20030 28022 20062
rect 15232 19992 15308 19998
rect 28021 19998 28022 20030
rect 28086 20030 28092 20062
rect 28696 20270 28702 20302
rect 28766 20302 28767 20334
rect 28968 20334 29044 20340
rect 28766 20270 28772 20302
rect 28696 20062 28772 20270
rect 28086 19998 28087 20030
rect 28021 19997 28087 19998
rect 28696 19998 28702 20062
rect 28766 19998 28772 20062
rect 28968 20270 28974 20334
rect 29038 20270 29044 20334
rect 28968 20062 29044 20270
rect 28968 20030 28974 20062
rect 28696 19992 28772 19998
rect 28973 19998 28974 20030
rect 29038 20030 29044 20062
rect 29240 20334 29316 20340
rect 29240 20270 29246 20334
rect 29310 20270 29316 20334
rect 29240 20062 29316 20270
rect 29240 20030 29246 20062
rect 29038 19998 29039 20030
rect 28973 19997 29039 19998
rect 29245 19998 29246 20030
rect 29310 20030 29316 20062
rect 29310 19998 29311 20030
rect 29245 19997 29311 19998
rect 14144 19926 14220 19932
rect 14144 19862 14150 19926
rect 14214 19862 14220 19926
rect 14557 19926 14623 19927
rect 14557 19894 14558 19926
rect 14144 19654 14220 19862
rect 14144 19622 14150 19654
rect 14149 19590 14150 19622
rect 14214 19622 14220 19654
rect 14552 19862 14558 19894
rect 14622 19894 14623 19926
rect 15096 19926 15172 19932
rect 14622 19862 14628 19894
rect 14552 19654 14628 19862
rect 14214 19590 14215 19622
rect 14149 19589 14215 19590
rect 14552 19590 14558 19654
rect 14622 19590 14628 19654
rect 15096 19862 15102 19926
rect 15166 19862 15172 19926
rect 15237 19926 15303 19927
rect 15237 19894 15238 19926
rect 15096 19654 15172 19862
rect 15096 19622 15102 19654
rect 14552 19584 14628 19590
rect 15101 19590 15102 19622
rect 15166 19622 15172 19654
rect 15232 19862 15238 19894
rect 15302 19894 15303 19926
rect 28293 19926 28359 19927
rect 28293 19894 28294 19926
rect 15302 19862 15308 19894
rect 15232 19654 15308 19862
rect 15166 19590 15167 19622
rect 15101 19589 15167 19590
rect 15232 19590 15238 19654
rect 15302 19590 15308 19654
rect 15232 19584 15308 19590
rect 28288 19862 28294 19894
rect 28358 19894 28359 19926
rect 28424 19926 28500 19932
rect 28358 19862 28364 19894
rect 28288 19654 28364 19862
rect 28288 19590 28294 19654
rect 28358 19590 28364 19654
rect 28424 19862 28430 19926
rect 28494 19862 28500 19926
rect 28837 19926 28903 19927
rect 28837 19894 28838 19926
rect 28424 19654 28500 19862
rect 28424 19622 28430 19654
rect 28288 19584 28364 19590
rect 28429 19590 28430 19622
rect 28494 19622 28500 19654
rect 28832 19862 28838 19894
rect 28902 19894 28903 19926
rect 29245 19926 29311 19927
rect 29245 19894 29246 19926
rect 28902 19862 28908 19894
rect 28832 19654 28908 19862
rect 28494 19590 28495 19622
rect 28429 19589 28495 19590
rect 28832 19590 28838 19654
rect 28902 19590 28908 19654
rect 28832 19584 28908 19590
rect 29240 19862 29246 19894
rect 29310 19894 29311 19926
rect 29310 19862 29316 19894
rect 29240 19654 29316 19862
rect 29240 19590 29246 19654
rect 29310 19590 29316 19654
rect 29240 19584 29316 19590
rect 14149 19518 14215 19519
rect 14149 19486 14150 19518
rect 14144 19454 14150 19486
rect 14214 19486 14215 19518
rect 14552 19518 14628 19524
rect 14214 19454 14220 19486
rect 14144 19246 14220 19454
rect 14144 19182 14150 19246
rect 14214 19182 14220 19246
rect 14552 19454 14558 19518
rect 14622 19454 14628 19518
rect 14552 19246 14628 19454
rect 14552 19214 14558 19246
rect 14144 19176 14220 19182
rect 14557 19182 14558 19214
rect 14622 19214 14628 19246
rect 14960 19518 15036 19524
rect 14960 19454 14966 19518
rect 15030 19454 15036 19518
rect 14960 19246 15036 19454
rect 14960 19214 14966 19246
rect 14622 19182 14623 19214
rect 14557 19181 14623 19182
rect 14965 19182 14966 19214
rect 15030 19214 15036 19246
rect 15232 19518 15308 19524
rect 15232 19454 15238 19518
rect 15302 19454 15308 19518
rect 28157 19518 28223 19519
rect 28157 19486 28158 19518
rect 15232 19246 15308 19454
rect 15232 19214 15238 19246
rect 15030 19182 15031 19214
rect 14965 19181 15031 19182
rect 15237 19182 15238 19214
rect 15302 19214 15308 19246
rect 28152 19454 28158 19486
rect 28222 19486 28223 19518
rect 28429 19518 28495 19519
rect 28429 19486 28430 19518
rect 28222 19454 28228 19486
rect 28152 19246 28228 19454
rect 15302 19182 15303 19214
rect 15237 19181 15303 19182
rect 28152 19182 28158 19246
rect 28222 19182 28228 19246
rect 28152 19176 28228 19182
rect 28424 19454 28430 19486
rect 28494 19486 28495 19518
rect 28832 19518 28908 19524
rect 28494 19454 28500 19486
rect 28424 19246 28500 19454
rect 28424 19182 28430 19246
rect 28494 19182 28500 19246
rect 28832 19454 28838 19518
rect 28902 19454 28908 19518
rect 28832 19246 28908 19454
rect 28832 19214 28838 19246
rect 28424 19176 28500 19182
rect 28837 19182 28838 19214
rect 28902 19214 28908 19246
rect 29240 19518 29316 19524
rect 29240 19454 29246 19518
rect 29310 19454 29316 19518
rect 29240 19246 29316 19454
rect 29240 19214 29246 19246
rect 28902 19182 28903 19214
rect 28837 19181 28903 19182
rect 29245 19182 29246 19214
rect 29310 19214 29316 19246
rect 29310 19182 29311 19214
rect 29245 19181 29311 19182
rect 14965 19110 15031 19111
rect 14965 19078 14966 19110
rect 14960 19046 14966 19078
rect 15030 19078 15031 19110
rect 15232 19110 15308 19116
rect 15030 19046 15036 19078
rect 14960 18838 15036 19046
rect 14960 18774 14966 18838
rect 15030 18774 15036 18838
rect 15232 19046 15238 19110
rect 15302 19046 15308 19110
rect 15232 18838 15308 19046
rect 28016 19110 28092 19116
rect 28016 19046 28022 19110
rect 28086 19046 28092 19110
rect 15232 18806 15238 18838
rect 14960 18768 15036 18774
rect 15237 18774 15238 18806
rect 15302 18806 15308 18838
rect 25160 18974 25236 18980
rect 25160 18910 25166 18974
rect 25230 18910 25236 18974
rect 15302 18774 15303 18806
rect 15237 18773 15303 18774
rect 15101 18702 15167 18703
rect 15101 18670 15102 18702
rect 12240 18502 12246 18566
rect 12310 18502 12316 18566
rect 12240 18496 12316 18502
rect 15096 18638 15102 18670
rect 15166 18670 15167 18702
rect 15373 18702 15439 18703
rect 15373 18670 15374 18702
rect 15166 18638 15172 18670
rect 15096 18430 15172 18638
rect 15096 18366 15102 18430
rect 15166 18366 15172 18430
rect 15096 18360 15172 18366
rect 15368 18638 15374 18670
rect 15438 18670 15439 18702
rect 25160 18702 25236 18910
rect 28016 18838 28092 19046
rect 28016 18806 28022 18838
rect 28021 18774 28022 18806
rect 28086 18806 28092 18838
rect 28424 19110 28500 19116
rect 28424 19046 28430 19110
rect 28494 19046 28500 19110
rect 28424 18838 28500 19046
rect 28424 18806 28430 18838
rect 28086 18774 28087 18806
rect 28021 18773 28087 18774
rect 28429 18774 28430 18806
rect 28494 18806 28500 18838
rect 28494 18774 28495 18806
rect 28429 18773 28495 18774
rect 25160 18670 25166 18702
rect 15438 18638 15444 18670
rect 15368 18430 15444 18638
rect 25165 18638 25166 18670
rect 25230 18670 25236 18702
rect 28152 18702 28228 18708
rect 25230 18638 25231 18670
rect 25165 18637 25231 18638
rect 28152 18638 28158 18702
rect 28222 18638 28228 18702
rect 28701 18702 28767 18703
rect 28701 18670 28702 18702
rect 15781 18566 15847 18567
rect 15781 18534 15782 18566
rect 15368 18366 15374 18430
rect 15438 18366 15444 18430
rect 15368 18360 15444 18366
rect 15776 18502 15782 18534
rect 15846 18534 15847 18566
rect 27880 18566 27956 18572
rect 15846 18502 15852 18534
rect 10472 17686 10478 17750
rect 10542 17686 10548 17750
rect 11832 18294 11908 18300
rect 11832 18230 11838 18294
rect 11902 18230 11908 18294
rect 11832 17750 11908 18230
rect 11832 17718 11838 17750
rect 10472 17680 10548 17686
rect 11837 17686 11838 17718
rect 11902 17718 11908 17750
rect 12240 18294 12316 18300
rect 12240 18230 12246 18294
rect 12310 18230 12316 18294
rect 12381 18294 12447 18295
rect 12381 18262 12382 18294
rect 11902 17686 11903 17718
rect 11837 17685 11903 17686
rect 12240 17478 12316 18230
rect 12376 18230 12382 18262
rect 12446 18262 12447 18294
rect 12517 18294 12583 18295
rect 12517 18262 12518 18294
rect 12446 18230 12452 18262
rect 12376 17750 12452 18230
rect 12376 17686 12382 17750
rect 12446 17686 12452 17750
rect 12376 17680 12452 17686
rect 12512 18230 12518 18262
rect 12582 18262 12583 18294
rect 12582 18230 12588 18262
rect 12512 17750 12588 18230
rect 14149 18022 14215 18023
rect 14149 17990 14150 18022
rect 12512 17686 12518 17750
rect 12582 17686 12588 17750
rect 12512 17680 12588 17686
rect 14144 17958 14150 17990
rect 14214 17990 14215 18022
rect 14688 18022 14764 18028
rect 14214 17958 14220 17990
rect 14144 17750 14220 17958
rect 14144 17686 14150 17750
rect 14214 17686 14220 17750
rect 14688 17958 14694 18022
rect 14758 17958 14764 18022
rect 14688 17750 14764 17958
rect 15776 18022 15852 18502
rect 27880 18502 27886 18566
rect 27950 18502 27956 18566
rect 18224 18430 18300 18436
rect 18224 18366 18230 18430
rect 18294 18366 18300 18430
rect 16189 18294 16255 18295
rect 16189 18262 16190 18294
rect 15776 17958 15782 18022
rect 15846 17958 15852 18022
rect 15776 17952 15852 17958
rect 16184 18230 16190 18262
rect 16254 18262 16255 18294
rect 16254 18230 16260 18262
rect 16184 18022 16260 18230
rect 18224 18158 18300 18366
rect 27613 18294 27679 18295
rect 27613 18262 27614 18294
rect 18224 18126 18230 18158
rect 18229 18094 18230 18126
rect 18294 18126 18300 18158
rect 27608 18230 27614 18262
rect 27678 18262 27679 18294
rect 27678 18230 27684 18262
rect 18294 18094 18295 18126
rect 18229 18093 18295 18094
rect 16184 17958 16190 18022
rect 16254 17958 16260 18022
rect 16184 17952 16260 17958
rect 26520 18022 26596 18028
rect 26520 17958 26526 18022
rect 26590 17958 26596 18022
rect 14688 17718 14694 17750
rect 14144 17680 14220 17686
rect 14693 17686 14694 17718
rect 14758 17718 14764 17750
rect 18365 17750 18431 17751
rect 18365 17718 18366 17750
rect 14758 17686 14759 17718
rect 14693 17685 14759 17686
rect 18360 17686 18366 17718
rect 18430 17718 18431 17750
rect 25296 17750 25372 17756
rect 18430 17686 18436 17718
rect 14144 17614 14220 17620
rect 14144 17550 14150 17614
rect 14214 17550 14220 17614
rect 14693 17614 14759 17615
rect 14693 17582 14694 17614
rect 12240 17446 12246 17478
rect 12245 17414 12246 17446
rect 12310 17446 12316 17478
rect 12648 17478 12724 17484
rect 12310 17414 12311 17446
rect 12245 17413 12311 17414
rect 12648 17414 12654 17478
rect 12718 17414 12724 17478
rect 12648 16118 12724 17414
rect 12648 16086 12654 16118
rect 12653 16054 12654 16086
rect 12718 16086 12724 16118
rect 13056 17478 13132 17484
rect 13056 17414 13062 17478
rect 13126 17414 13132 17478
rect 13056 16118 13132 17414
rect 14144 17342 14220 17550
rect 14144 17310 14150 17342
rect 14149 17278 14150 17310
rect 14214 17310 14220 17342
rect 14688 17550 14694 17582
rect 14758 17582 14759 17614
rect 14758 17550 14764 17582
rect 14688 17342 14764 17550
rect 18360 17478 18436 17686
rect 18360 17414 18366 17478
rect 18430 17414 18436 17478
rect 25296 17686 25302 17750
rect 25366 17686 25372 17750
rect 26520 17750 26596 17958
rect 27608 18022 27684 18230
rect 27608 17958 27614 18022
rect 27678 17958 27684 18022
rect 27880 18022 27956 18502
rect 28152 18430 28228 18638
rect 28152 18398 28158 18430
rect 28157 18366 28158 18398
rect 28222 18398 28228 18430
rect 28696 18638 28702 18670
rect 28766 18670 28767 18702
rect 28766 18638 28772 18670
rect 28696 18430 28772 18638
rect 28222 18366 28223 18398
rect 28157 18365 28223 18366
rect 28696 18366 28702 18430
rect 28766 18366 28772 18430
rect 28696 18360 28772 18366
rect 30469 18294 30535 18295
rect 30469 18262 30470 18294
rect 30464 18230 30470 18262
rect 30534 18262 30535 18294
rect 31149 18294 31215 18295
rect 31149 18262 31150 18294
rect 30534 18230 30540 18262
rect 27880 17990 27886 18022
rect 27608 17952 27684 17958
rect 27885 17958 27886 17990
rect 27950 17990 27956 18022
rect 28973 18022 29039 18023
rect 28973 17990 28974 18022
rect 27950 17958 27951 17990
rect 27885 17957 27951 17958
rect 28968 17958 28974 17990
rect 29038 17990 29039 18022
rect 29240 18022 29316 18028
rect 29038 17958 29044 17990
rect 26520 17718 26526 17750
rect 25296 17478 25372 17686
rect 26525 17686 26526 17718
rect 26590 17718 26596 17750
rect 28968 17750 29044 17958
rect 26590 17686 26591 17718
rect 26525 17685 26591 17686
rect 28968 17686 28974 17750
rect 29038 17686 29044 17750
rect 29240 17958 29246 18022
rect 29310 17958 29316 18022
rect 29240 17750 29316 17958
rect 29240 17718 29246 17750
rect 28968 17680 29044 17686
rect 29245 17686 29246 17718
rect 29310 17718 29316 17750
rect 30464 17750 30540 18230
rect 29310 17686 29311 17718
rect 29245 17685 29311 17686
rect 30464 17686 30470 17750
rect 30534 17686 30540 17750
rect 30464 17680 30540 17686
rect 31144 18230 31150 18262
rect 31214 18262 31215 18294
rect 31693 18294 31759 18295
rect 31693 18262 31694 18294
rect 31214 18230 31220 18262
rect 31144 17750 31220 18230
rect 31144 17686 31150 17750
rect 31214 17686 31220 17750
rect 31144 17680 31220 17686
rect 31688 18230 31694 18262
rect 31758 18262 31759 18294
rect 31758 18230 31764 18262
rect 31688 17750 31764 18230
rect 31688 17686 31694 17750
rect 31758 17686 31764 17750
rect 31688 17680 31764 17686
rect 39848 17750 39924 17756
rect 39848 17686 39854 17750
rect 39918 17686 39924 17750
rect 28973 17614 29039 17615
rect 28973 17582 28974 17614
rect 25296 17446 25302 17478
rect 18360 17408 18436 17414
rect 25301 17414 25302 17446
rect 25366 17446 25372 17478
rect 28968 17550 28974 17582
rect 29038 17582 29039 17614
rect 29245 17614 29311 17615
rect 29245 17582 29246 17614
rect 29038 17550 29044 17582
rect 25366 17414 25367 17446
rect 25301 17413 25367 17414
rect 14214 17278 14215 17310
rect 14149 17277 14215 17278
rect 14688 17278 14694 17342
rect 14758 17278 14764 17342
rect 14688 17272 14764 17278
rect 18360 17342 18436 17348
rect 18360 17278 18366 17342
rect 18430 17278 18436 17342
rect 25301 17342 25367 17343
rect 25301 17310 25302 17342
rect 14285 17206 14351 17207
rect 14285 17174 14286 17206
rect 14280 17142 14286 17174
rect 14350 17174 14351 17206
rect 14688 17206 14764 17212
rect 14350 17142 14356 17174
rect 14280 16934 14356 17142
rect 14280 16870 14286 16934
rect 14350 16870 14356 16934
rect 14688 17142 14694 17206
rect 14758 17142 14764 17206
rect 15101 17206 15167 17207
rect 15101 17174 15102 17206
rect 14688 16934 14764 17142
rect 14688 16902 14694 16934
rect 14280 16864 14356 16870
rect 14693 16870 14694 16902
rect 14758 16902 14764 16934
rect 15096 17142 15102 17174
rect 15166 17174 15167 17206
rect 15232 17206 15308 17212
rect 15166 17142 15172 17174
rect 15096 16934 15172 17142
rect 14758 16870 14759 16902
rect 14693 16869 14759 16870
rect 15096 16870 15102 16934
rect 15166 16870 15172 16934
rect 15232 17142 15238 17206
rect 15302 17142 15308 17206
rect 15232 16934 15308 17142
rect 18360 17070 18436 17278
rect 18360 17038 18366 17070
rect 18365 17006 18366 17038
rect 18430 17038 18436 17070
rect 25296 17278 25302 17310
rect 25366 17310 25367 17342
rect 28968 17342 29044 17550
rect 25366 17278 25372 17310
rect 25296 17070 25372 17278
rect 28968 17278 28974 17342
rect 29038 17278 29044 17342
rect 28968 17272 29044 17278
rect 29240 17550 29246 17582
rect 29310 17582 29311 17614
rect 29310 17550 29316 17582
rect 29240 17342 29316 17550
rect 30469 17478 30535 17479
rect 30469 17446 30470 17478
rect 29240 17278 29246 17342
rect 29310 17278 29316 17342
rect 29240 17272 29316 17278
rect 30464 17414 30470 17446
rect 30534 17446 30535 17478
rect 30872 17478 30948 17484
rect 30534 17414 30540 17446
rect 18430 17006 18431 17038
rect 18365 17005 18431 17006
rect 25296 17006 25302 17070
rect 25366 17006 25372 17070
rect 25296 17000 25372 17006
rect 28152 17206 28228 17212
rect 28152 17142 28158 17206
rect 28222 17142 28228 17206
rect 15232 16902 15238 16934
rect 15096 16864 15172 16870
rect 15237 16870 15238 16902
rect 15302 16902 15308 16934
rect 28152 16934 28228 17142
rect 28152 16902 28158 16934
rect 15302 16870 15303 16902
rect 15237 16869 15303 16870
rect 28157 16870 28158 16902
rect 28222 16902 28228 16934
rect 28696 17206 28772 17212
rect 28696 17142 28702 17206
rect 28766 17142 28772 17206
rect 28973 17206 29039 17207
rect 28973 17174 28974 17206
rect 28696 16934 28772 17142
rect 28696 16902 28702 16934
rect 28222 16870 28223 16902
rect 28157 16869 28223 16870
rect 28701 16870 28702 16902
rect 28766 16902 28772 16934
rect 28968 17142 28974 17174
rect 29038 17174 29039 17206
rect 29240 17206 29316 17212
rect 29038 17142 29044 17174
rect 28968 16934 29044 17142
rect 28766 16870 28767 16902
rect 28701 16869 28767 16870
rect 28968 16870 28974 16934
rect 29038 16870 29044 16934
rect 29240 17142 29246 17206
rect 29310 17142 29316 17206
rect 29240 16934 29316 17142
rect 29240 16902 29246 16934
rect 28968 16864 29044 16870
rect 29245 16870 29246 16902
rect 29310 16902 29316 16934
rect 29310 16870 29311 16902
rect 29245 16869 29311 16870
rect 14144 16798 14220 16804
rect 14144 16734 14150 16798
rect 14214 16734 14220 16798
rect 14557 16798 14623 16799
rect 14557 16766 14558 16798
rect 14144 16526 14220 16734
rect 14144 16494 14150 16526
rect 14149 16462 14150 16494
rect 14214 16494 14220 16526
rect 14552 16734 14558 16766
rect 14622 16766 14623 16798
rect 15101 16798 15167 16799
rect 15101 16766 15102 16798
rect 14622 16734 14628 16766
rect 14552 16526 14628 16734
rect 14214 16462 14215 16494
rect 14149 16461 14215 16462
rect 14552 16462 14558 16526
rect 14622 16462 14628 16526
rect 14552 16456 14628 16462
rect 15096 16734 15102 16766
rect 15166 16766 15167 16798
rect 15504 16798 15580 16804
rect 15166 16734 15172 16766
rect 15096 16526 15172 16734
rect 15096 16462 15102 16526
rect 15166 16462 15172 16526
rect 15504 16734 15510 16798
rect 15574 16734 15580 16798
rect 28157 16798 28223 16799
rect 28157 16766 28158 16798
rect 15504 16526 15580 16734
rect 15504 16494 15510 16526
rect 15096 16456 15172 16462
rect 15509 16462 15510 16494
rect 15574 16494 15580 16526
rect 28152 16734 28158 16766
rect 28222 16766 28223 16798
rect 28565 16798 28631 16799
rect 28565 16766 28566 16798
rect 28222 16734 28228 16766
rect 28152 16526 28228 16734
rect 15574 16462 15575 16494
rect 15509 16461 15575 16462
rect 28152 16462 28158 16526
rect 28222 16462 28228 16526
rect 28152 16456 28228 16462
rect 28560 16734 28566 16766
rect 28630 16766 28631 16798
rect 28973 16798 29039 16799
rect 28973 16766 28974 16798
rect 28630 16734 28636 16766
rect 28560 16526 28636 16734
rect 28560 16462 28566 16526
rect 28630 16462 28636 16526
rect 28560 16456 28636 16462
rect 28968 16734 28974 16766
rect 29038 16766 29039 16798
rect 29240 16798 29316 16804
rect 29038 16734 29044 16766
rect 28968 16526 29044 16734
rect 28968 16462 28974 16526
rect 29038 16462 29044 16526
rect 29240 16734 29246 16798
rect 29310 16734 29316 16798
rect 29240 16526 29316 16734
rect 29240 16494 29246 16526
rect 28968 16456 29044 16462
rect 29245 16462 29246 16494
rect 29310 16494 29316 16526
rect 29310 16462 29311 16494
rect 29245 16461 29311 16462
rect 14285 16390 14351 16391
rect 14285 16358 14286 16390
rect 13056 16086 13062 16118
rect 12718 16054 12719 16086
rect 12653 16053 12719 16054
rect 13061 16054 13062 16086
rect 13126 16086 13132 16118
rect 14280 16326 14286 16358
rect 14350 16358 14351 16390
rect 14688 16390 14764 16396
rect 14350 16326 14356 16358
rect 14280 16118 14356 16326
rect 13126 16054 13127 16086
rect 13061 16053 13127 16054
rect 14280 16054 14286 16118
rect 14350 16054 14356 16118
rect 14688 16326 14694 16390
rect 14758 16326 14764 16390
rect 14688 16118 14764 16326
rect 14688 16086 14694 16118
rect 14280 16048 14356 16054
rect 14693 16054 14694 16086
rect 14758 16086 14764 16118
rect 15096 16390 15172 16396
rect 15096 16326 15102 16390
rect 15166 16326 15172 16390
rect 15509 16390 15575 16391
rect 15509 16358 15510 16390
rect 15096 16118 15172 16326
rect 15096 16086 15102 16118
rect 14758 16054 14759 16086
rect 14693 16053 14759 16054
rect 15101 16054 15102 16086
rect 15166 16086 15172 16118
rect 15504 16326 15510 16358
rect 15574 16358 15575 16390
rect 28293 16390 28359 16391
rect 28293 16358 28294 16390
rect 15574 16326 15580 16358
rect 15504 16118 15580 16326
rect 15166 16054 15167 16086
rect 15101 16053 15167 16054
rect 15504 16054 15510 16118
rect 15574 16054 15580 16118
rect 15504 16048 15580 16054
rect 28288 16326 28294 16358
rect 28358 16358 28359 16390
rect 28560 16390 28636 16396
rect 28358 16326 28364 16358
rect 28288 16118 28364 16326
rect 28288 16054 28294 16118
rect 28358 16054 28364 16118
rect 28560 16326 28566 16390
rect 28630 16326 28636 16390
rect 28560 16118 28636 16326
rect 28560 16086 28566 16118
rect 28288 16048 28364 16054
rect 28565 16054 28566 16086
rect 28630 16086 28636 16118
rect 28968 16390 29044 16396
rect 28968 16326 28974 16390
rect 29038 16326 29044 16390
rect 28968 16118 29044 16326
rect 28968 16086 28974 16118
rect 28630 16054 28631 16086
rect 28565 16053 28631 16054
rect 28973 16054 28974 16086
rect 29038 16086 29044 16118
rect 29240 16390 29316 16396
rect 29240 16326 29246 16390
rect 29310 16326 29316 16390
rect 29240 16118 29316 16326
rect 29240 16086 29246 16118
rect 29038 16054 29039 16086
rect 28973 16053 29039 16054
rect 29245 16054 29246 16086
rect 29310 16086 29316 16118
rect 30464 16118 30540 17414
rect 29310 16054 29311 16086
rect 29245 16053 29311 16054
rect 30464 16054 30470 16118
rect 30534 16054 30540 16118
rect 30872 17414 30878 17478
rect 30942 17414 30948 17478
rect 30872 16118 30948 17414
rect 30872 16086 30878 16118
rect 30464 16048 30540 16054
rect 30877 16054 30878 16086
rect 30942 16086 30948 16118
rect 30942 16054 30943 16086
rect 30877 16053 30943 16054
rect 3808 15374 3814 15438
rect 3878 15374 3884 15438
rect 3808 15368 3884 15374
rect 11968 15982 12044 15988
rect 11968 15918 11974 15982
rect 12038 15918 12044 15982
rect 3405 15302 3471 15303
rect 3405 15270 3406 15302
rect 3400 15238 3406 15270
rect 3470 15270 3471 15302
rect 11968 15302 12044 15918
rect 11968 15270 11974 15302
rect 3470 15238 3476 15270
rect 2640 12938 2706 12939
rect 2640 12874 2641 12938
rect 2705 12874 2706 12938
rect 2640 12873 2706 12874
rect 3400 12582 3476 15238
rect 11973 15238 11974 15270
rect 12038 15270 12044 15302
rect 12240 15982 12316 15988
rect 12240 15918 12246 15982
rect 12310 15918 12316 15982
rect 12789 15982 12855 15983
rect 12789 15950 12790 15982
rect 12240 15302 12316 15918
rect 12784 15918 12790 15950
rect 12854 15950 12855 15982
rect 14280 15982 14356 15988
rect 12854 15918 12860 15950
rect 12784 15710 12860 15918
rect 12784 15646 12790 15710
rect 12854 15646 12860 15710
rect 14280 15918 14286 15982
rect 14350 15918 14356 15982
rect 14693 15982 14759 15983
rect 14693 15950 14694 15982
rect 14280 15710 14356 15918
rect 14280 15678 14286 15710
rect 12784 15640 12860 15646
rect 14285 15646 14286 15678
rect 14350 15678 14356 15710
rect 14688 15918 14694 15950
rect 14758 15950 14759 15982
rect 14965 15982 15031 15983
rect 14965 15950 14966 15982
rect 14758 15918 14764 15950
rect 14688 15710 14764 15918
rect 14350 15646 14351 15678
rect 14285 15645 14351 15646
rect 14688 15646 14694 15710
rect 14758 15646 14764 15710
rect 14688 15640 14764 15646
rect 14960 15918 14966 15950
rect 15030 15950 15031 15982
rect 15504 15982 15580 15988
rect 15030 15918 15036 15950
rect 14960 15710 15036 15918
rect 14960 15646 14966 15710
rect 15030 15646 15036 15710
rect 15504 15918 15510 15982
rect 15574 15918 15580 15982
rect 28157 15982 28223 15983
rect 28157 15950 28158 15982
rect 15504 15710 15580 15918
rect 15504 15678 15510 15710
rect 14960 15640 15036 15646
rect 15509 15646 15510 15678
rect 15574 15678 15580 15710
rect 28152 15918 28158 15950
rect 28222 15950 28223 15982
rect 28560 15982 28636 15988
rect 28222 15918 28228 15950
rect 28152 15710 28228 15918
rect 15574 15646 15575 15678
rect 15509 15645 15575 15646
rect 28152 15646 28158 15710
rect 28222 15646 28228 15710
rect 28560 15918 28566 15982
rect 28630 15918 28636 15982
rect 28973 15982 29039 15983
rect 28973 15950 28974 15982
rect 28560 15710 28636 15918
rect 28560 15678 28566 15710
rect 28152 15640 28228 15646
rect 28565 15646 28566 15678
rect 28630 15678 28636 15710
rect 28968 15918 28974 15950
rect 29038 15950 29039 15982
rect 29376 15982 29452 15988
rect 29038 15918 29044 15950
rect 28968 15710 29044 15918
rect 28630 15646 28631 15678
rect 28565 15645 28631 15646
rect 28968 15646 28974 15710
rect 29038 15646 29044 15710
rect 29376 15918 29382 15982
rect 29446 15918 29452 15982
rect 29376 15710 29452 15918
rect 29376 15678 29382 15710
rect 28968 15640 29044 15646
rect 29381 15646 29382 15678
rect 29446 15678 29452 15710
rect 31008 15982 31084 15988
rect 31008 15918 31014 15982
rect 31078 15918 31084 15982
rect 29446 15646 29447 15678
rect 29381 15645 29447 15646
rect 14149 15574 14215 15575
rect 14149 15542 14150 15574
rect 12240 15270 12246 15302
rect 12038 15238 12039 15270
rect 11973 15237 12039 15238
rect 12245 15238 12246 15270
rect 12310 15270 12316 15302
rect 14144 15510 14150 15542
rect 14214 15542 14215 15574
rect 14688 15574 14764 15580
rect 14214 15510 14220 15542
rect 14144 15302 14220 15510
rect 12310 15238 12311 15270
rect 12245 15237 12311 15238
rect 14144 15238 14150 15302
rect 14214 15238 14220 15302
rect 14688 15510 14694 15574
rect 14758 15510 14764 15574
rect 14965 15574 15031 15575
rect 14965 15542 14966 15574
rect 14688 15302 14764 15510
rect 14688 15270 14694 15302
rect 14144 15232 14220 15238
rect 14693 15238 14694 15270
rect 14758 15270 14764 15302
rect 14960 15510 14966 15542
rect 15030 15542 15031 15574
rect 15237 15574 15303 15575
rect 15237 15542 15238 15574
rect 15030 15510 15036 15542
rect 14960 15302 15036 15510
rect 14758 15238 14759 15270
rect 14693 15237 14759 15238
rect 14960 15238 14966 15302
rect 15030 15238 15036 15302
rect 14960 15232 15036 15238
rect 15232 15510 15238 15542
rect 15302 15542 15303 15574
rect 28016 15574 28092 15580
rect 15302 15510 15308 15542
rect 15232 15302 15308 15510
rect 15232 15238 15238 15302
rect 15302 15238 15308 15302
rect 28016 15510 28022 15574
rect 28086 15510 28092 15574
rect 28565 15574 28631 15575
rect 28565 15542 28566 15574
rect 28016 15302 28092 15510
rect 28016 15270 28022 15302
rect 15232 15232 15308 15238
rect 28021 15238 28022 15270
rect 28086 15270 28092 15302
rect 28560 15510 28566 15542
rect 28630 15542 28631 15574
rect 28968 15574 29044 15580
rect 28630 15510 28636 15542
rect 28560 15302 28636 15510
rect 28086 15238 28087 15270
rect 28021 15237 28087 15238
rect 28560 15238 28566 15302
rect 28630 15238 28636 15302
rect 28968 15510 28974 15574
rect 29038 15510 29044 15574
rect 29245 15574 29311 15575
rect 29245 15542 29246 15574
rect 28968 15302 29044 15510
rect 28968 15270 28974 15302
rect 28560 15232 28636 15238
rect 28973 15238 28974 15270
rect 29038 15270 29044 15302
rect 29240 15510 29246 15542
rect 29310 15542 29311 15574
rect 29310 15510 29316 15542
rect 29240 15302 29316 15510
rect 29038 15238 29039 15270
rect 28973 15237 29039 15238
rect 29240 15238 29246 15302
rect 29310 15238 29316 15302
rect 31008 15302 31084 15918
rect 31008 15270 31014 15302
rect 29240 15232 29316 15238
rect 31013 15238 31014 15270
rect 31078 15270 31084 15302
rect 31280 15982 31356 15988
rect 31280 15918 31286 15982
rect 31350 15918 31356 15982
rect 31280 15302 31356 15918
rect 31280 15270 31286 15302
rect 31078 15238 31079 15270
rect 31013 15237 31079 15238
rect 31285 15238 31286 15270
rect 31350 15270 31356 15302
rect 31350 15238 31351 15270
rect 31285 15237 31351 15238
rect 10472 15166 10548 15172
rect 10472 15102 10478 15166
rect 10542 15102 10548 15166
rect 10472 14078 10548 15102
rect 10472 14046 10478 14078
rect 10477 14014 10478 14046
rect 10542 14046 10548 14078
rect 10880 15166 10956 15172
rect 10880 15102 10886 15166
rect 10950 15102 10956 15166
rect 12109 15166 12175 15167
rect 12109 15134 12110 15166
rect 10542 14014 10543 14046
rect 10477 14013 10543 14014
rect 9525 13806 9591 13807
rect 9525 13774 9526 13806
rect 3400 12518 3406 12582
rect 3470 12518 3476 12582
rect 3400 12512 3476 12518
rect 9520 13742 9526 13774
rect 9590 13774 9591 13806
rect 9590 13742 9596 13774
rect 4085 12446 4151 12447
rect 4085 12414 4086 12446
rect 952 12246 1230 12310
rect 1294 12246 1300 12310
rect 952 10406 1300 12246
rect 4080 12382 4086 12414
rect 4150 12414 4151 12446
rect 9384 12446 9460 12452
rect 4150 12382 4156 12414
rect 3264 11086 3340 11092
rect 3264 11022 3270 11086
rect 3334 11022 3340 11086
rect 3264 10542 3340 11022
rect 3264 10510 3270 10542
rect 3269 10478 3270 10510
rect 3334 10510 3340 10542
rect 3334 10478 3335 10510
rect 3269 10477 3335 10478
rect 952 10342 1230 10406
rect 1294 10342 1300 10406
rect 952 8910 1300 10342
rect 4080 9726 4156 12382
rect 4080 9662 4086 9726
rect 4150 9662 4156 9726
rect 9384 12382 9390 12446
rect 9454 12382 9460 12446
rect 9384 9726 9460 12382
rect 9520 11222 9596 13742
rect 10880 12582 10956 15102
rect 12104 15102 12110 15134
rect 12174 15134 12175 15166
rect 12512 15166 12588 15172
rect 12174 15102 12180 15134
rect 12104 14894 12180 15102
rect 12104 14830 12110 14894
rect 12174 14830 12180 14894
rect 12512 15102 12518 15166
rect 12582 15102 12588 15166
rect 15373 15166 15439 15167
rect 15373 15134 15374 15166
rect 12512 14894 12588 15102
rect 12512 14862 12518 14894
rect 12104 14824 12180 14830
rect 12517 14830 12518 14862
rect 12582 14862 12588 14894
rect 15368 15102 15374 15134
rect 15438 15134 15439 15166
rect 32781 15166 32847 15167
rect 32781 15134 32782 15166
rect 15438 15102 15444 15134
rect 12582 14830 12583 14862
rect 12517 14829 12583 14830
rect 15368 14758 15444 15102
rect 32776 15102 32782 15134
rect 32846 15134 32847 15166
rect 34685 15166 34751 15167
rect 34685 15134 34686 15166
rect 32846 15102 32852 15134
rect 15368 14694 15374 14758
rect 15438 14694 15444 14758
rect 15368 14688 15444 14694
rect 18224 15030 18300 15036
rect 18224 14966 18230 15030
rect 18294 14966 18300 15030
rect 17685 14622 17751 14623
rect 17685 14590 17686 14622
rect 17680 14558 17686 14590
rect 17750 14590 17751 14622
rect 18224 14622 18300 14966
rect 19589 14758 19655 14759
rect 19589 14726 19590 14758
rect 18224 14590 18230 14622
rect 17750 14558 17756 14590
rect 17680 14350 17756 14558
rect 18229 14558 18230 14590
rect 18294 14590 18300 14622
rect 19584 14694 19590 14726
rect 19654 14726 19655 14758
rect 25160 14758 25236 14764
rect 19654 14694 19660 14726
rect 18294 14558 18295 14590
rect 18229 14557 18295 14558
rect 17680 14286 17686 14350
rect 17750 14286 17756 14350
rect 17680 14280 17756 14286
rect 19045 14214 19111 14215
rect 19045 14182 19046 14214
rect 19040 14150 19046 14182
rect 19110 14182 19111 14214
rect 19110 14150 19116 14182
rect 19040 13806 19116 14150
rect 19040 13742 19046 13806
rect 19110 13742 19116 13806
rect 19040 13736 19116 13742
rect 10880 12550 10886 12582
rect 10885 12518 10886 12550
rect 10950 12550 10956 12582
rect 19584 12582 19660 14694
rect 25160 14694 25166 14758
rect 25230 14694 25236 14758
rect 20808 14214 20884 14220
rect 20808 14150 20814 14214
rect 20878 14150 20884 14214
rect 21493 14214 21559 14215
rect 21493 14182 21494 14214
rect 20808 13806 20884 14150
rect 20808 13774 20814 13806
rect 20813 13742 20814 13774
rect 20878 13774 20884 13806
rect 21488 14150 21494 14182
rect 21558 14182 21559 14214
rect 22032 14214 22108 14220
rect 21558 14150 21564 14182
rect 21488 13806 21564 14150
rect 20878 13742 20879 13774
rect 20813 13741 20879 13742
rect 21488 13742 21494 13806
rect 21558 13742 21564 13806
rect 22032 14150 22038 14214
rect 22102 14150 22108 14214
rect 22717 14214 22783 14215
rect 22717 14182 22718 14214
rect 22032 13806 22108 14150
rect 22032 13774 22038 13806
rect 21488 13736 21564 13742
rect 22037 13742 22038 13774
rect 22102 13774 22108 13806
rect 22712 14150 22718 14182
rect 22782 14182 22783 14214
rect 23125 14214 23191 14215
rect 23125 14182 23126 14214
rect 22782 14150 22788 14182
rect 22712 13806 22788 14150
rect 22102 13742 22103 13774
rect 22037 13741 22103 13742
rect 22712 13742 22718 13806
rect 22782 13742 22788 13806
rect 22712 13736 22788 13742
rect 23120 14150 23126 14182
rect 23190 14182 23191 14214
rect 23256 14214 23332 14220
rect 23190 14150 23196 14182
rect 23120 13806 23196 14150
rect 23120 13742 23126 13806
rect 23190 13742 23196 13806
rect 23256 14150 23262 14214
rect 23326 14150 23332 14214
rect 23805 14214 23871 14215
rect 23805 14182 23806 14214
rect 23256 13806 23332 14150
rect 23256 13774 23262 13806
rect 23120 13736 23196 13742
rect 23261 13742 23262 13774
rect 23326 13774 23332 13806
rect 23800 14150 23806 14182
rect 23870 14182 23871 14214
rect 23941 14214 24007 14215
rect 23941 14182 23942 14214
rect 23870 14150 23876 14182
rect 23800 13806 23876 14150
rect 23326 13742 23327 13774
rect 23261 13741 23327 13742
rect 23800 13742 23806 13806
rect 23870 13742 23876 13806
rect 23800 13736 23876 13742
rect 23936 14150 23942 14182
rect 24006 14182 24007 14214
rect 24006 14150 24012 14182
rect 23936 13806 24012 14150
rect 23936 13742 23942 13806
rect 24006 13742 24012 13806
rect 23936 13736 24012 13742
rect 22581 13670 22647 13671
rect 22581 13638 22582 13670
rect 22576 13606 22582 13638
rect 22646 13638 22647 13670
rect 22646 13606 22652 13638
rect 10950 12518 10951 12550
rect 10885 12517 10951 12518
rect 19584 12518 19590 12582
rect 19654 12518 19660 12582
rect 20133 12582 20199 12583
rect 20133 12550 20134 12582
rect 19584 12512 19660 12518
rect 20128 12518 20134 12550
rect 20198 12550 20199 12582
rect 20198 12518 20204 12550
rect 9520 11158 9526 11222
rect 9590 11158 9596 11222
rect 9520 11152 9596 11158
rect 9525 11086 9591 11087
rect 9525 11054 9526 11086
rect 9384 9694 9390 9726
rect 4080 9656 4156 9662
rect 9389 9662 9390 9694
rect 9454 9694 9460 9726
rect 9520 11022 9526 11054
rect 9590 11054 9591 11086
rect 9590 11022 9596 11054
rect 9454 9662 9455 9694
rect 9389 9661 9455 9662
rect 952 8846 1230 8910
rect 1294 8846 1300 8910
rect 952 7142 1300 8846
rect 9384 9590 9460 9596
rect 9384 9526 9390 9590
rect 9454 9526 9460 9590
rect 3269 8774 3335 8775
rect 3269 8742 3270 8774
rect 3264 8710 3270 8742
rect 3334 8742 3335 8774
rect 3334 8710 3340 8742
rect 3264 8366 3340 8710
rect 3264 8302 3270 8366
rect 3334 8302 3340 8366
rect 3264 8296 3340 8302
rect 952 7078 1230 7142
rect 1294 7078 1300 7142
rect 952 5374 1300 7078
rect 9384 7006 9460 9526
rect 9520 8366 9596 11022
rect 19992 10950 20068 10956
rect 19992 10886 19998 10950
rect 20062 10886 20068 10950
rect 19725 10814 19791 10815
rect 19725 10782 19726 10814
rect 19720 10750 19726 10782
rect 19790 10782 19791 10814
rect 19790 10750 19796 10782
rect 9520 8302 9526 8366
rect 9590 8302 9596 8366
rect 9520 8296 9596 8302
rect 19040 8774 19116 8780
rect 19040 8710 19046 8774
rect 19110 8710 19116 8774
rect 9384 6974 9390 7006
rect 9389 6942 9390 6974
rect 9454 6974 9460 7006
rect 9520 8230 9596 8236
rect 9520 8166 9526 8230
rect 9590 8166 9596 8230
rect 9454 6942 9455 6974
rect 9389 6941 9455 6942
rect 9520 6876 9596 8166
rect 19040 7006 19116 8710
rect 19312 8502 19388 8508
rect 19312 8438 19318 8502
rect 19382 8438 19388 8502
rect 19312 8094 19388 8438
rect 19312 8062 19318 8094
rect 19317 8030 19318 8062
rect 19382 8062 19388 8094
rect 19382 8030 19383 8062
rect 19317 8029 19383 8030
rect 19040 6974 19046 7006
rect 19045 6942 19046 6974
rect 19110 6974 19116 7006
rect 19110 6942 19111 6974
rect 19045 6941 19111 6942
rect 9384 6800 9596 6876
rect 9384 5510 9460 6800
rect 9525 6734 9591 6735
rect 9525 6702 9526 6734
rect 9384 5478 9390 5510
rect 9389 5446 9390 5478
rect 9454 5478 9460 5510
rect 9520 6670 9526 6702
rect 9590 6702 9591 6734
rect 9590 6670 9596 6702
rect 9454 5446 9455 5478
rect 9389 5445 9455 5446
rect 952 5310 1230 5374
rect 1294 5310 1300 5374
rect 9253 5374 9319 5375
rect 9253 5342 9254 5374
rect 952 3878 1300 5310
rect 952 3814 1230 3878
rect 1294 3814 1300 3878
rect 952 1294 1300 3814
rect 9248 5310 9254 5342
rect 9318 5342 9319 5374
rect 9318 5310 9324 5342
rect 5989 3198 6055 3199
rect 5989 3166 5990 3198
rect 5984 3134 5990 3166
rect 6054 3166 6055 3198
rect 6054 3134 6060 3166
rect 2045 2110 2111 2111
rect 2045 2078 2046 2110
rect 2040 2046 2046 2078
rect 2110 2078 2111 2110
rect 2110 2046 2116 2078
rect 2040 1838 2116 2046
rect 2040 1774 2046 1838
rect 2110 1774 2116 1838
rect 2040 1768 2116 1774
rect 2181 1702 2247 1703
rect 2181 1670 2182 1702
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 1300 1294
rect 952 1158 1300 1230
rect 2176 1638 2182 1670
rect 2246 1670 2247 1702
rect 3813 1702 3879 1703
rect 3813 1670 3814 1702
rect 2246 1638 2252 1670
rect 2176 1294 2252 1638
rect 2176 1230 2182 1294
rect 2246 1230 2252 1294
rect 2176 1224 2252 1230
rect 3808 1638 3814 1670
rect 3878 1670 3879 1702
rect 5445 1702 5511 1703
rect 5445 1670 5446 1702
rect 3878 1638 3884 1670
rect 3808 1294 3884 1638
rect 3808 1230 3814 1294
rect 3878 1230 3884 1294
rect 3808 1224 3884 1230
rect 5440 1638 5446 1670
rect 5510 1670 5511 1702
rect 5510 1638 5516 1670
rect 5440 1294 5516 1638
rect 5440 1230 5446 1294
rect 5510 1230 5516 1294
rect 5440 1224 5516 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 1300 1158
rect 952 1022 1300 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 1300 1022
rect 952 952 1300 958
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 620 614
rect 272 478 620 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 620 478
rect 272 342 620 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 620 342
rect 272 272 620 278
rect 5984 0 6060 3134
rect 9248 2654 9324 5310
rect 9520 4150 9596 6670
rect 9520 4086 9526 4150
rect 9590 4086 9596 4150
rect 9520 4080 9596 4086
rect 9248 2590 9254 2654
rect 9318 2590 9324 2654
rect 9248 2584 9324 2590
rect 9384 4014 9460 4020
rect 9384 3950 9390 4014
rect 9454 3950 9460 4014
rect 9384 1838 9460 3950
rect 10749 3198 10815 3199
rect 10749 3166 10750 3198
rect 10744 3134 10750 3166
rect 10814 3166 10815 3198
rect 12109 3198 12175 3199
rect 12109 3166 12110 3198
rect 10814 3134 10820 3166
rect 9525 2518 9591 2519
rect 9525 2486 9526 2518
rect 9384 1806 9390 1838
rect 9389 1774 9390 1806
rect 9454 1806 9460 1838
rect 9520 2454 9526 2486
rect 9590 2486 9591 2518
rect 9590 2454 9596 2486
rect 9454 1774 9455 1806
rect 9389 1773 9455 1774
rect 7077 1702 7143 1703
rect 7077 1670 7078 1702
rect 7072 1638 7078 1670
rect 7142 1670 7143 1702
rect 8709 1702 8775 1703
rect 8709 1670 8710 1702
rect 7142 1638 7148 1670
rect 7072 1294 7148 1638
rect 7072 1230 7078 1294
rect 7142 1230 7148 1294
rect 7072 1224 7148 1230
rect 8704 1638 8710 1670
rect 8774 1670 8775 1702
rect 8774 1638 8780 1670
rect 8704 1294 8780 1638
rect 8704 1230 8710 1294
rect 8774 1230 8780 1294
rect 8704 1224 8780 1230
rect 9520 614 9596 2454
rect 10341 1702 10407 1703
rect 10341 1670 10342 1702
rect 10336 1638 10342 1670
rect 10406 1670 10407 1702
rect 10406 1638 10412 1670
rect 10336 1294 10412 1638
rect 10336 1230 10342 1294
rect 10406 1230 10412 1294
rect 10336 1224 10412 1230
rect 9520 550 9526 614
rect 9590 550 9596 614
rect 9520 544 9596 550
rect 10744 0 10820 3134
rect 12104 3134 12110 3166
rect 12174 3166 12175 3198
rect 13197 3198 13263 3199
rect 13197 3166 13198 3198
rect 12174 3134 12180 3166
rect 12104 0 12180 3134
rect 13192 3134 13198 3166
rect 13262 3166 13263 3198
rect 14421 3198 14487 3199
rect 14421 3166 14422 3198
rect 13262 3134 13268 3166
rect 12245 1702 12311 1703
rect 12245 1670 12246 1702
rect 12240 1638 12246 1670
rect 12310 1670 12311 1702
rect 12310 1638 12316 1670
rect 12240 1294 12316 1638
rect 12240 1230 12246 1294
rect 12310 1230 12316 1294
rect 12240 1224 12316 1230
rect 13192 0 13268 3134
rect 14416 3134 14422 3166
rect 14486 3166 14487 3198
rect 15509 3198 15575 3199
rect 15509 3166 15510 3198
rect 14486 3134 14492 3166
rect 13741 1702 13807 1703
rect 13741 1670 13742 1702
rect 13736 1638 13742 1670
rect 13806 1670 13807 1702
rect 13806 1638 13812 1670
rect 13736 1294 13812 1638
rect 13736 1230 13742 1294
rect 13806 1230 13812 1294
rect 13736 1224 13812 1230
rect 14416 0 14492 3134
rect 15504 3134 15510 3166
rect 15574 3166 15575 3198
rect 16733 3198 16799 3199
rect 16733 3166 16734 3198
rect 15574 3134 15580 3166
rect 15373 1702 15439 1703
rect 15373 1670 15374 1702
rect 15368 1638 15374 1670
rect 15438 1670 15439 1702
rect 15438 1638 15444 1670
rect 15368 1294 15444 1638
rect 15368 1230 15374 1294
rect 15438 1230 15444 1294
rect 15368 1224 15444 1230
rect 15504 0 15580 3134
rect 16728 3134 16734 3166
rect 16798 3166 16799 3198
rect 17957 3198 18023 3199
rect 17957 3166 17958 3198
rect 16798 3134 16804 3166
rect 16728 0 16804 3134
rect 17952 3134 17958 3166
rect 18022 3166 18023 3198
rect 19045 3198 19111 3199
rect 19045 3166 19046 3198
rect 18022 3134 18028 3166
rect 17277 1702 17343 1703
rect 17277 1670 17278 1702
rect 17272 1638 17278 1670
rect 17342 1670 17343 1702
rect 17342 1638 17348 1670
rect 17272 1294 17348 1638
rect 17272 1230 17278 1294
rect 17342 1230 17348 1294
rect 17272 1224 17348 1230
rect 17952 0 18028 3134
rect 19040 3134 19046 3166
rect 19110 3166 19111 3198
rect 19110 3134 19116 3166
rect 18773 1702 18839 1703
rect 18773 1670 18774 1702
rect 18768 1638 18774 1670
rect 18838 1670 18839 1702
rect 18838 1638 18844 1670
rect 18768 1294 18844 1638
rect 18768 1230 18774 1294
rect 18838 1230 18844 1294
rect 18768 1224 18844 1230
rect 19040 0 19116 3134
rect 19720 0 19796 10750
rect 19992 9590 20068 10886
rect 20128 10678 20204 12518
rect 22576 11902 22652 13606
rect 25160 12582 25236 14694
rect 32776 13534 32852 15102
rect 34680 15102 34686 15134
rect 34750 15134 34751 15166
rect 39848 15166 39924 17686
rect 39848 15134 39854 15166
rect 34750 15102 34756 15134
rect 34680 14894 34756 15102
rect 39853 15102 39854 15134
rect 39918 15134 39924 15166
rect 39918 15102 39919 15134
rect 39853 15101 39919 15102
rect 34680 14830 34686 14894
rect 34750 14830 34756 14894
rect 34680 14824 34756 14830
rect 40120 14894 40196 14900
rect 40120 14830 40126 14894
rect 40190 14830 40196 14894
rect 34685 14758 34751 14759
rect 34685 14726 34686 14758
rect 32776 13470 32782 13534
rect 32846 13470 32852 13534
rect 32776 13464 32852 13470
rect 34680 14694 34686 14726
rect 34750 14726 34751 14758
rect 34750 14694 34756 14726
rect 25160 12550 25166 12582
rect 25165 12518 25166 12550
rect 25230 12550 25236 12582
rect 25230 12518 25231 12550
rect 25165 12517 25231 12518
rect 34680 12174 34756 14694
rect 34680 12110 34686 12174
rect 34750 12110 34756 12174
rect 34680 12104 34756 12110
rect 34816 13398 34892 13404
rect 34816 13334 34822 13398
rect 34886 13334 34892 13398
rect 22576 11838 22582 11902
rect 22646 11838 22652 11902
rect 22576 11832 22652 11838
rect 34680 11902 34756 11908
rect 34680 11838 34686 11902
rect 34750 11838 34756 11902
rect 20264 11766 20340 11772
rect 20264 11702 20270 11766
rect 20334 11702 20340 11766
rect 20264 11086 20340 11702
rect 20264 11054 20270 11086
rect 20269 11022 20270 11054
rect 20334 11054 20340 11086
rect 20334 11022 20335 11054
rect 20269 11021 20335 11022
rect 20949 10814 21015 10815
rect 20949 10782 20950 10814
rect 20128 10614 20134 10678
rect 20198 10614 20204 10678
rect 20128 10608 20204 10614
rect 20944 10750 20950 10782
rect 21014 10782 21015 10814
rect 22445 10814 22511 10815
rect 22445 10782 22446 10814
rect 21014 10750 21020 10782
rect 20128 10542 20204 10548
rect 20128 10478 20134 10542
rect 20198 10478 20204 10542
rect 20269 10542 20335 10543
rect 20269 10510 20270 10542
rect 20128 9998 20204 10478
rect 20128 9966 20134 9998
rect 20133 9934 20134 9966
rect 20198 9966 20204 9998
rect 20264 10478 20270 10510
rect 20334 10510 20335 10542
rect 20334 10478 20340 10510
rect 20198 9934 20199 9966
rect 20133 9933 20199 9934
rect 19992 9558 19998 9590
rect 19997 9526 19998 9558
rect 20062 9558 20068 9590
rect 20128 9726 20204 9732
rect 20128 9662 20134 9726
rect 20198 9662 20204 9726
rect 20062 9526 20063 9558
rect 19997 9525 20063 9526
rect 20128 9182 20204 9662
rect 20128 9150 20134 9182
rect 20133 9118 20134 9150
rect 20198 9150 20204 9182
rect 20198 9118 20199 9150
rect 20133 9117 20199 9118
rect 20264 3340 20340 10478
rect 20813 9726 20879 9727
rect 20813 9694 20814 9726
rect 20808 9662 20814 9694
rect 20878 9694 20879 9726
rect 20878 9662 20884 9694
rect 20677 9318 20743 9319
rect 20677 9286 20678 9318
rect 20672 9254 20678 9286
rect 20742 9286 20743 9318
rect 20742 9254 20748 9286
rect 20672 8502 20748 9254
rect 20808 9182 20884 9662
rect 20808 9118 20814 9182
rect 20878 9118 20884 9182
rect 20808 9112 20884 9118
rect 20672 8438 20678 8502
rect 20742 8438 20748 8502
rect 20672 8432 20748 8438
rect 20264 3264 20476 3340
rect 20269 3198 20335 3199
rect 20269 3166 20270 3198
rect 20264 3134 20270 3166
rect 20334 3166 20335 3198
rect 20334 3134 20340 3166
rect 20264 0 20340 3134
rect 20400 0 20476 3264
rect 20677 1702 20743 1703
rect 20677 1670 20678 1702
rect 20672 1638 20678 1670
rect 20742 1670 20743 1702
rect 20742 1638 20748 1670
rect 20672 1294 20748 1638
rect 20672 1230 20678 1294
rect 20742 1230 20748 1294
rect 20672 1224 20748 1230
rect 20944 0 21020 10750
rect 22440 10750 22446 10782
rect 22510 10782 22511 10814
rect 23669 10814 23735 10815
rect 23669 10782 23670 10814
rect 22510 10750 22516 10782
rect 21493 10542 21559 10543
rect 21493 10510 21494 10542
rect 21488 10478 21494 10510
rect 21558 10510 21559 10542
rect 21629 10542 21695 10543
rect 21629 10510 21630 10542
rect 21558 10478 21564 10510
rect 21488 10134 21564 10478
rect 21488 10070 21494 10134
rect 21558 10070 21564 10134
rect 21488 10064 21564 10070
rect 21624 10478 21630 10510
rect 21694 10510 21695 10542
rect 22168 10542 22244 10548
rect 21694 10478 21700 10510
rect 21357 3198 21423 3199
rect 21357 3166 21358 3198
rect 21352 3134 21358 3166
rect 21422 3166 21423 3198
rect 21422 3134 21428 3166
rect 21352 0 21428 3134
rect 21624 0 21700 10478
rect 22168 10478 22174 10542
rect 22238 10478 22244 10542
rect 22168 9998 22244 10478
rect 22168 9966 22174 9998
rect 22173 9934 22174 9966
rect 22238 9966 22244 9998
rect 22238 9934 22239 9966
rect 22173 9933 22239 9934
rect 22309 1702 22375 1703
rect 22309 1670 22310 1702
rect 22304 1638 22310 1670
rect 22374 1670 22375 1702
rect 22374 1638 22380 1670
rect 22304 1294 22380 1638
rect 22304 1230 22310 1294
rect 22374 1230 22380 1294
rect 22304 1224 22380 1230
rect 22440 0 22516 10750
rect 23664 10750 23670 10782
rect 23734 10782 23735 10814
rect 23734 10750 23740 10782
rect 22712 10542 22788 10548
rect 22712 10478 22718 10542
rect 22782 10478 22788 10542
rect 22853 10542 22919 10543
rect 22853 10510 22854 10542
rect 22712 9998 22788 10478
rect 22712 9966 22718 9998
rect 22717 9934 22718 9966
rect 22782 9966 22788 9998
rect 22848 10478 22854 10510
rect 22918 10510 22919 10542
rect 23392 10542 23468 10548
rect 22918 10478 22924 10510
rect 22782 9934 22783 9966
rect 22717 9933 22783 9934
rect 22581 3198 22647 3199
rect 22581 3166 22582 3198
rect 22576 3134 22582 3166
rect 22646 3166 22647 3198
rect 22646 3134 22652 3166
rect 22576 0 22652 3134
rect 22848 0 22924 10478
rect 23392 10478 23398 10542
rect 23462 10478 23468 10542
rect 23392 10270 23468 10478
rect 23392 10238 23398 10270
rect 23397 10206 23398 10238
rect 23462 10238 23468 10270
rect 23462 10206 23463 10238
rect 23397 10205 23463 10206
rect 23261 9726 23327 9727
rect 23261 9694 23262 9726
rect 23256 9662 23262 9694
rect 23326 9694 23327 9726
rect 23326 9662 23332 9694
rect 23256 9182 23332 9662
rect 23256 9118 23262 9182
rect 23326 9118 23332 9182
rect 23256 9112 23332 9118
rect 23533 1702 23599 1703
rect 23533 1670 23534 1702
rect 23528 1638 23534 1670
rect 23598 1670 23599 1702
rect 23598 1638 23604 1670
rect 23528 1294 23604 1638
rect 23528 1230 23534 1294
rect 23598 1230 23604 1294
rect 23528 1224 23604 1230
rect 23664 0 23740 10750
rect 23936 10542 24012 10548
rect 23936 10478 23942 10542
rect 24006 10478 24012 10542
rect 24077 10542 24143 10543
rect 24077 10510 24078 10542
rect 23936 9998 24012 10478
rect 23936 9966 23942 9998
rect 23941 9934 23942 9966
rect 24006 9966 24012 9998
rect 24072 10478 24078 10510
rect 24142 10510 24143 10542
rect 24142 10478 24148 10510
rect 24006 9934 24007 9966
rect 23941 9933 24007 9934
rect 23805 3198 23871 3199
rect 23805 3166 23806 3198
rect 23800 3134 23806 3166
rect 23870 3166 23871 3198
rect 23870 3134 23876 3166
rect 23800 0 23876 3134
rect 24072 0 24148 10478
rect 34680 9318 34756 11838
rect 34816 10678 34892 13334
rect 40120 12310 40196 14830
rect 40795 12864 40855 23033
rect 42160 22238 42508 23806
rect 42160 22174 42166 22238
rect 42230 22174 42508 22238
rect 42160 20470 42508 22174
rect 42160 20406 42166 20470
rect 42230 20406 42508 20470
rect 41621 19246 41687 19247
rect 41621 19214 41622 19246
rect 41616 19182 41622 19214
rect 41686 19214 41687 19246
rect 41686 19182 41692 19214
rect 41616 18974 41692 19182
rect 41616 18910 41622 18974
rect 41686 18910 41692 18974
rect 41616 18904 41692 18910
rect 42160 18974 42508 20406
rect 42160 18910 42166 18974
rect 42230 18910 42508 18974
rect 41616 17206 41692 17212
rect 41616 17142 41622 17206
rect 41686 17142 41692 17206
rect 41616 16526 41692 17142
rect 41616 16494 41622 16526
rect 41621 16462 41622 16494
rect 41686 16494 41692 16526
rect 42160 17206 42508 18910
rect 42160 17142 42166 17206
rect 42230 17142 42508 17206
rect 41686 16462 41687 16494
rect 41621 16461 41687 16462
rect 42160 15438 42508 17142
rect 42160 15374 42166 15438
rect 42230 15374 42508 15438
rect 42160 13806 42508 15374
rect 42160 13742 42166 13806
rect 42230 13742 42508 13806
rect 40792 12863 40858 12864
rect 40792 12799 40793 12863
rect 40857 12799 40858 12863
rect 40792 12798 40858 12799
rect 40120 12278 40126 12310
rect 40125 12246 40126 12278
rect 40190 12278 40196 12310
rect 42160 12310 42508 13742
rect 40190 12246 40191 12278
rect 40125 12245 40191 12246
rect 42160 12246 42166 12310
rect 42230 12246 42508 12310
rect 34816 10646 34822 10678
rect 34821 10614 34822 10646
rect 34886 10646 34892 10678
rect 34886 10614 34887 10646
rect 34821 10613 34887 10614
rect 34680 9286 34686 9318
rect 34685 9254 34686 9286
rect 34750 9286 34756 9318
rect 42160 10406 42508 12246
rect 42160 10342 42166 10406
rect 42230 10342 42508 10406
rect 34750 9254 34751 9286
rect 34685 9253 34751 9254
rect 24485 8774 24551 8775
rect 24485 8742 24486 8774
rect 24480 8710 24486 8742
rect 24550 8742 24551 8774
rect 42160 8774 42508 10342
rect 24550 8710 24556 8742
rect 24349 8502 24415 8503
rect 24349 8470 24350 8502
rect 24344 8438 24350 8470
rect 24414 8470 24415 8502
rect 24414 8438 24420 8470
rect 24344 8094 24420 8438
rect 24344 8030 24350 8094
rect 24414 8030 24420 8094
rect 24344 8024 24420 8030
rect 24480 7006 24556 8710
rect 24480 6942 24486 7006
rect 24550 6942 24556 7006
rect 24480 6936 24556 6942
rect 42160 8710 42166 8774
rect 42230 8710 42508 8774
rect 42160 7142 42508 8710
rect 42160 7078 42166 7142
rect 42230 7078 42508 7142
rect 42160 5374 42508 7078
rect 42160 5310 42166 5374
rect 42230 5310 42508 5374
rect 42160 3878 42508 5310
rect 42160 3814 42166 3878
rect 42230 3814 42508 3878
rect 42160 2110 42508 3814
rect 42160 2046 42166 2110
rect 42230 2046 42508 2110
rect 25437 1702 25503 1703
rect 25437 1670 25438 1702
rect 25432 1638 25438 1670
rect 25502 1670 25503 1702
rect 27341 1702 27407 1703
rect 27341 1670 27342 1702
rect 25502 1638 25508 1670
rect 25432 1294 25508 1638
rect 25432 1230 25438 1294
rect 25502 1230 25508 1294
rect 25432 1224 25508 1230
rect 27336 1638 27342 1670
rect 27406 1670 27407 1702
rect 28973 1702 29039 1703
rect 28973 1670 28974 1702
rect 27406 1638 27412 1670
rect 27336 1294 27412 1638
rect 27336 1230 27342 1294
rect 27406 1230 27412 1294
rect 27336 1224 27412 1230
rect 28968 1638 28974 1670
rect 29038 1670 29039 1702
rect 30605 1702 30671 1703
rect 30605 1670 30606 1702
rect 29038 1638 29044 1670
rect 28968 1294 29044 1638
rect 28968 1230 28974 1294
rect 29038 1230 29044 1294
rect 28968 1224 29044 1230
rect 30600 1638 30606 1670
rect 30670 1670 30671 1702
rect 32237 1702 32303 1703
rect 32237 1670 32238 1702
rect 30670 1638 30676 1670
rect 30600 1294 30676 1638
rect 30600 1230 30606 1294
rect 30670 1230 30676 1294
rect 30600 1224 30676 1230
rect 32232 1638 32238 1670
rect 32302 1670 32303 1702
rect 34005 1702 34071 1703
rect 34005 1670 34006 1702
rect 32302 1638 32308 1670
rect 32232 1294 32308 1638
rect 32232 1230 32238 1294
rect 32302 1230 32308 1294
rect 32232 1224 32308 1230
rect 34000 1638 34006 1670
rect 34070 1670 34071 1702
rect 35637 1702 35703 1703
rect 35637 1670 35638 1702
rect 34070 1638 34076 1670
rect 34000 1294 34076 1638
rect 34000 1230 34006 1294
rect 34070 1230 34076 1294
rect 34000 1224 34076 1230
rect 35632 1638 35638 1670
rect 35702 1670 35703 1702
rect 37405 1702 37471 1703
rect 37405 1670 37406 1702
rect 35702 1638 35708 1670
rect 35632 1294 35708 1638
rect 35632 1230 35638 1294
rect 35702 1230 35708 1294
rect 35632 1224 35708 1230
rect 37400 1638 37406 1670
rect 37470 1670 37471 1702
rect 39037 1702 39103 1703
rect 39037 1670 39038 1702
rect 37470 1638 37476 1670
rect 37400 1294 37476 1638
rect 37400 1230 37406 1294
rect 37470 1230 37476 1294
rect 37400 1224 37476 1230
rect 39032 1638 39038 1670
rect 39102 1670 39103 1702
rect 40805 1702 40871 1703
rect 40805 1670 40806 1702
rect 39102 1638 39108 1670
rect 39032 1294 39108 1638
rect 39032 1230 39038 1294
rect 39102 1230 39108 1294
rect 39032 1224 39108 1230
rect 40800 1638 40806 1670
rect 40870 1670 40871 1702
rect 40870 1638 40876 1670
rect 40800 1294 40876 1638
rect 40800 1230 40806 1294
rect 40870 1230 40876 1294
rect 40800 1224 40876 1230
rect 42160 1294 42508 2046
rect 42160 1230 42166 1294
rect 42230 1230 42302 1294
rect 42366 1230 42438 1294
rect 42502 1230 42508 1294
rect 42160 1158 42508 1230
rect 42160 1094 42166 1158
rect 42230 1094 42302 1158
rect 42366 1094 42438 1158
rect 42502 1094 42508 1158
rect 42160 1022 42508 1094
rect 42160 958 42166 1022
rect 42230 958 42302 1022
rect 42366 958 42438 1022
rect 42502 958 42508 1022
rect 42160 952 42508 958
rect 42840 30534 43188 32510
rect 42840 30470 42846 30534
rect 42910 30470 43188 30534
rect 42840 23462 43188 30470
rect 42840 23398 42846 23462
rect 42910 23398 43188 23462
rect 42840 17886 43188 23398
rect 42840 17822 42846 17886
rect 42910 17822 43188 17886
rect 42840 614 43188 17822
rect 42840 550 42846 614
rect 42910 550 42982 614
rect 43046 550 43118 614
rect 43182 550 43188 614
rect 42840 478 43188 550
rect 42840 414 42846 478
rect 42910 414 42982 478
rect 43046 414 43118 478
rect 43182 414 43188 478
rect 42840 342 43188 414
rect 42840 278 42846 342
rect 42910 278 42982 342
rect 43046 278 43118 342
rect 43182 278 43188 342
rect 42840 272 43188 278
use contact_30  contact_30_0
timestamp 1634918361
transform 1 0 42840 0 1 30469
box 0 0 1 1
use contact_30  contact_30_1
timestamp 1634918361
transform 1 0 40120 0 1 14829
box 0 0 1 1
use contact_30  contact_30_2
timestamp 1634918361
transform 1 0 40120 0 1 12245
box 0 0 1 1
use contact_30  contact_30_3
timestamp 1634918361
transform 1 0 42840 0 1 17821
box 0 0 1 1
use contact_30  contact_30_4
timestamp 1634918361
transform 1 0 42840 0 1 23397
box 0 0 1 1
use contact_30  contact_30_5
timestamp 1634918361
transform 1 0 40120 0 1 20677
box 0 0 1 1
use contact_30  contact_30_6
timestamp 1634918361
transform 1 0 40120 0 1 23397
box 0 0 1 1
use contact_30  contact_30_7
timestamp 1634918361
transform 1 0 39848 0 1 17685
box 0 0 1 1
use contact_30  contact_30_8
timestamp 1634918361
transform 1 0 39848 0 1 15101
box 0 0 1 1
use contact_30  contact_30_9
timestamp 1634918361
transform 1 0 34680 0 1 11837
box 0 0 1 1
use contact_30  contact_30_10
timestamp 1634918361
transform 1 0 34680 0 1 9253
box 0 0 1 1
use contact_30  contact_30_11
timestamp 1634918361
transform 1 0 34680 0 1 12109
box 0 0 1 1
use contact_30  contact_30_12
timestamp 1634918361
transform 1 0 34680 0 1 14693
box 0 0 1 1
use contact_30  contact_30_13
timestamp 1634918361
transform 1 0 34272 0 1 32509
box 0 0 1 1
use contact_30  contact_30_14
timestamp 1634918361
transform 1 0 34272 0 1 30605
box 0 0 1 1
use contact_30  contact_30_15
timestamp 1634918361
transform 1 0 34000 0 1 27749
box 0 0 1 1
use contact_30  contact_30_16
timestamp 1634918361
transform 1 0 34000 0 1 30469
box 0 0 1 1
use contact_30  contact_30_17
timestamp 1634918361
transform 1 0 34408 0 1 27613
box 0 0 1 1
use contact_30  contact_30_18
timestamp 1634918361
transform 1 0 34408 0 1 24893
box 0 0 1 1
use contact_30  contact_30_19
timestamp 1634918361
transform 1 0 34272 0 1 24757
box 0 0 1 1
use contact_30  contact_30_20
timestamp 1634918361
transform 1 0 34272 0 1 22173
box 0 0 1 1
use contact_30  contact_30_21
timestamp 1634918361
transform 1 0 34680 0 1 14829
box 0 0 1 1
use contact_30  contact_30_22
timestamp 1634918361
transform 1 0 34680 0 1 15101
box 0 0 1 1
use contact_30  contact_30_23
timestamp 1634918361
transform 1 0 31688 0 1 17685
box 0 0 1 1
use contact_30  contact_30_24
timestamp 1634918361
transform 1 0 31688 0 1 18229
box 0 0 1 1
use contact_30  contact_30_25
timestamp 1634918361
transform 1 0 30872 0 1 17413
box 0 0 1 1
use contact_30  contact_30_26
timestamp 1634918361
transform 1 0 30872 0 1 16053
box 0 0 1 1
use contact_30  contact_30_27
timestamp 1634918361
transform 1 0 31008 0 1 15917
box 0 0 1 1
use contact_30  contact_30_28
timestamp 1634918361
transform 1 0 31008 0 1 15237
box 0 0 1 1
use contact_30  contact_30_29
timestamp 1634918361
transform 1 0 29376 0 1 20677
box 0 0 1 1
use contact_30  contact_30_30
timestamp 1634918361
transform 1 0 29376 0 1 20405
box 0 0 1 1
use contact_30  contact_30_31
timestamp 1634918361
transform 1 0 29240 0 1 17141
box 0 0 1 1
use contact_30  contact_30_32
timestamp 1634918361
transform 1 0 29240 0 1 16869
box 0 0 1 1
use contact_30  contact_30_33
timestamp 1634918361
transform 1 0 29240 0 1 19453
box 0 0 1 1
use contact_30  contact_30_34
timestamp 1634918361
transform 1 0 29240 0 1 19181
box 0 0 1 1
use contact_30  contact_30_35
timestamp 1634918361
transform 1 0 29240 0 1 19589
box 0 0 1 1
use contact_30  contact_30_36
timestamp 1634918361
transform 1 0 29240 0 1 19861
box 0 0 1 1
use contact_30  contact_30_37
timestamp 1634918361
transform 1 0 29240 0 1 20269
box 0 0 1 1
use contact_30  contact_30_38
timestamp 1634918361
transform 1 0 29240 0 1 19997
box 0 0 1 1
use contact_30  contact_30_39
timestamp 1634918361
transform 1 0 29240 0 1 16733
box 0 0 1 1
use contact_30  contact_30_40
timestamp 1634918361
transform 1 0 29240 0 1 16461
box 0 0 1 1
use contact_30  contact_30_41
timestamp 1634918361
transform 1 0 29240 0 1 16325
box 0 0 1 1
use contact_30  contact_30_42
timestamp 1634918361
transform 1 0 29240 0 1 16053
box 0 0 1 1
use contact_30  contact_30_43
timestamp 1634918361
transform 1 0 29240 0 1 15237
box 0 0 1 1
use contact_30  contact_30_44
timestamp 1634918361
transform 1 0 29240 0 1 15509
box 0 0 1 1
use contact_30  contact_30_45
timestamp 1634918361
transform 1 0 29376 0 1 15917
box 0 0 1 1
use contact_30  contact_30_46
timestamp 1634918361
transform 1 0 29376 0 1 15645
box 0 0 1 1
use contact_30  contact_30_47
timestamp 1634918361
transform 1 0 29240 0 1 17277
box 0 0 1 1
use contact_30  contact_30_48
timestamp 1634918361
transform 1 0 29240 0 1 17549
box 0 0 1 1
use contact_30  contact_30_49
timestamp 1634918361
transform 1 0 29240 0 1 17957
box 0 0 1 1
use contact_30  contact_30_50
timestamp 1634918361
transform 1 0 29240 0 1 17685
box 0 0 1 1
use contact_30  contact_30_51
timestamp 1634918361
transform 1 0 28696 0 1 20677
box 0 0 1 1
use contact_30  contact_30_52
timestamp 1634918361
transform 1 0 28696 0 1 20405
box 0 0 1 1
use contact_30  contact_30_53
timestamp 1634918361
transform 1 0 28696 0 1 19997
box 0 0 1 1
use contact_30  contact_30_54
timestamp 1634918361
transform 1 0 28696 0 1 20269
box 0 0 1 1
use contact_30  contact_30_55
timestamp 1634918361
transform 1 0 28560 0 1 16325
box 0 0 1 1
use contact_30  contact_30_56
timestamp 1634918361
transform 1 0 28560 0 1 16053
box 0 0 1 1
use contact_30  contact_30_57
timestamp 1634918361
transform 1 0 28696 0 1 17141
box 0 0 1 1
use contact_30  contact_30_58
timestamp 1634918361
transform 1 0 28696 0 1 16869
box 0 0 1 1
use contact_30  contact_30_59
timestamp 1634918361
transform 1 0 28560 0 1 16461
box 0 0 1 1
use contact_30  contact_30_60
timestamp 1634918361
transform 1 0 28560 0 1 16733
box 0 0 1 1
use contact_30  contact_30_61
timestamp 1634918361
transform 1 0 28424 0 1 19861
box 0 0 1 1
use contact_30  contact_30_62
timestamp 1634918361
transform 1 0 28424 0 1 19589
box 0 0 1 1
use contact_30  contact_30_63
timestamp 1634918361
transform 1 0 28424 0 1 19181
box 0 0 1 1
use contact_30  contact_30_64
timestamp 1634918361
transform 1 0 28424 0 1 19453
box 0 0 1 1
use contact_30  contact_30_65
timestamp 1634918361
transform 1 0 28560 0 1 15237
box 0 0 1 1
use contact_30  contact_30_66
timestamp 1634918361
transform 1 0 28560 0 1 15509
box 0 0 1 1
use contact_30  contact_30_67
timestamp 1634918361
transform 1 0 28560 0 1 15917
box 0 0 1 1
use contact_30  contact_30_68
timestamp 1634918361
transform 1 0 28560 0 1 15645
box 0 0 1 1
use contact_30  contact_30_69
timestamp 1634918361
transform 1 0 28696 0 1 18365
box 0 0 1 1
use contact_30  contact_30_70
timestamp 1634918361
transform 1 0 28696 0 1 18637
box 0 0 1 1
use contact_30  contact_30_71
timestamp 1634918361
transform 1 0 28424 0 1 19045
box 0 0 1 1
use contact_30  contact_30_72
timestamp 1634918361
transform 1 0 28424 0 1 18773
box 0 0 1 1
use contact_30  contact_30_73
timestamp 1634918361
transform 1 0 27880 0 1 18501
box 0 0 1 1
use contact_30  contact_30_74
timestamp 1634918361
transform 1 0 27880 0 1 17957
box 0 0 1 1
use contact_30  contact_30_75
timestamp 1634918361
transform 1 0 27608 0 1 17957
box 0 0 1 1
use contact_30  contact_30_76
timestamp 1634918361
transform 1 0 27608 0 1 18229
box 0 0 1 1
use contact_30  contact_30_77
timestamp 1634918361
transform 1 0 26520 0 1 17957
box 0 0 1 1
use contact_30  contact_30_78
timestamp 1634918361
transform 1 0 26520 0 1 17685
box 0 0 1 1
use contact_30  contact_30_79
timestamp 1634918361
transform 1 0 25296 0 1 17685
box 0 0 1 1
use contact_30  contact_30_80
timestamp 1634918361
transform 1 0 25296 0 1 17413
box 0 0 1 1
use contact_30  contact_30_81
timestamp 1634918361
transform 1 0 25296 0 1 17005
box 0 0 1 1
use contact_30  contact_30_82
timestamp 1634918361
transform 1 0 25296 0 1 17277
box 0 0 1 1
use contact_30  contact_30_83
timestamp 1634918361
transform 1 0 25160 0 1 18909
box 0 0 1 1
use contact_30  contact_30_84
timestamp 1634918361
transform 1 0 25160 0 1 18637
box 0 0 1 1
use contact_30  contact_30_85
timestamp 1634918361
transform 1 0 24480 0 1 6941
box 0 0 1 1
use contact_30  contact_30_86
timestamp 1634918361
transform 1 0 24480 0 1 8709
box 0 0 1 1
use contact_30  contact_30_87
timestamp 1634918361
transform 1 0 23936 0 1 10477
box 0 0 1 1
use contact_30  contact_30_88
timestamp 1634918361
transform 1 0 23936 0 1 9933
box 0 0 1 1
use contact_30  contact_30_89
timestamp 1634918361
transform 1 0 25160 0 1 14693
box 0 0 1 1
use contact_30  contact_30_90
timestamp 1634918361
transform 1 0 25160 0 1 12517
box 0 0 1 1
use contact_30  contact_30_91
timestamp 1634918361
transform 1 0 23936 0 1 25165
box 0 0 1 1
use contact_30  contact_30_92
timestamp 1634918361
transform 1 0 23936 0 1 23397
box 0 0 1 1
use contact_30  contact_30_93
timestamp 1634918361
transform 1 0 23256 0 1 9117
box 0 0 1 1
use contact_30  contact_30_94
timestamp 1634918361
transform 1 0 23256 0 1 9661
box 0 0 1 1
use contact_30  contact_30_95
timestamp 1634918361
transform 1 0 23392 0 1 25437
box 0 0 1 1
use contact_30  contact_30_96
timestamp 1634918361
transform 1 0 23392 0 1 25709
box 0 0 1 1
use contact_30  contact_30_97
timestamp 1634918361
transform 1 0 22712 0 1 25709
box 0 0 1 1
use contact_30  contact_30_98
timestamp 1634918361
transform 1 0 22712 0 1 25437
box 0 0 1 1
use contact_30  contact_30_99
timestamp 1634918361
transform 1 0 23392 0 1 10477
box 0 0 1 1
use contact_30  contact_30_100
timestamp 1634918361
transform 1 0 23392 0 1 10205
box 0 0 1 1
use contact_30  contact_30_101
timestamp 1634918361
transform 1 0 22712 0 1 10477
box 0 0 1 1
use contact_30  contact_30_102
timestamp 1634918361
transform 1 0 22712 0 1 9933
box 0 0 1 1
use contact_30  contact_30_103
timestamp 1634918361
transform 1 0 22168 0 1 10477
box 0 0 1 1
use contact_30  contact_30_104
timestamp 1634918361
transform 1 0 22168 0 1 9933
box 0 0 1 1
use contact_30  contact_30_105
timestamp 1634918361
transform 1 0 22168 0 1 25437
box 0 0 1 1
use contact_30  contact_30_106
timestamp 1634918361
transform 1 0 22168 0 1 25709
box 0 0 1 1
use contact_30  contact_30_107
timestamp 1634918361
transform 1 0 21488 0 1 25709
box 0 0 1 1
use contact_30  contact_30_108
timestamp 1634918361
transform 1 0 21488 0 1 25437
box 0 0 1 1
use contact_30  contact_30_109
timestamp 1634918361
transform 1 0 21488 0 1 10069
box 0 0 1 1
use contact_30  contact_30_110
timestamp 1634918361
transform 1 0 21488 0 1 10477
box 0 0 1 1
use contact_30  contact_30_111
timestamp 1634918361
transform 1 0 20808 0 1 9117
box 0 0 1 1
use contact_30  contact_30_112
timestamp 1634918361
transform 1 0 20808 0 1 9661
box 0 0 1 1
use contact_30  contact_30_113
timestamp 1634918361
transform 1 0 20944 0 1 25437
box 0 0 1 1
use contact_30  contact_30_114
timestamp 1634918361
transform 1 0 20944 0 1 25709
box 0 0 1 1
use contact_30  contact_30_115
timestamp 1634918361
transform 1 0 20128 0 1 25709
box 0 0 1 1
use contact_30  contact_30_116
timestamp 1634918361
transform 1 0 20128 0 1 25437
box 0 0 1 1
use contact_30  contact_30_117
timestamp 1634918361
transform 1 0 20128 0 1 10477
box 0 0 1 1
use contact_30  contact_30_118
timestamp 1634918361
transform 1 0 20128 0 1 9933
box 0 0 1 1
use contact_30  contact_30_119
timestamp 1634918361
transform 1 0 20128 0 1 10613
box 0 0 1 1
use contact_30  contact_30_120
timestamp 1634918361
transform 1 0 20128 0 1 12517
box 0 0 1 1
use contact_30  contact_30_121
timestamp 1634918361
transform 1 0 20128 0 1 9661
box 0 0 1 1
use contact_30  contact_30_122
timestamp 1634918361
transform 1 0 20128 0 1 9117
box 0 0 1 1
use contact_30  contact_30_123
timestamp 1634918361
transform 1 0 19584 0 1 12517
box 0 0 1 1
use contact_30  contact_30_124
timestamp 1634918361
transform 1 0 19584 0 1 14693
box 0 0 1 1
use contact_30  contact_30_125
timestamp 1634918361
transform 1 0 18360 0 1 17413
box 0 0 1 1
use contact_30  contact_30_126
timestamp 1634918361
transform 1 0 18360 0 1 17685
box 0 0 1 1
use contact_30  contact_30_127
timestamp 1634918361
transform 1 0 18224 0 1 18365
box 0 0 1 1
use contact_30  contact_30_128
timestamp 1634918361
transform 1 0 18224 0 1 18093
box 0 0 1 1
use contact_30  contact_30_129
timestamp 1634918361
transform 1 0 18360 0 1 17277
box 0 0 1 1
use contact_30  contact_30_130
timestamp 1634918361
transform 1 0 18360 0 1 17005
box 0 0 1 1
use contact_30  contact_30_131
timestamp 1634918361
transform 1 0 18224 0 1 14965
box 0 0 1 1
use contact_30  contact_30_132
timestamp 1634918361
transform 1 0 18224 0 1 14557
box 0 0 1 1
use contact_30  contact_30_133
timestamp 1634918361
transform 1 0 19720 0 1 23397
box 0 0 1 1
use contact_30  contact_30_134
timestamp 1634918361
transform 1 0 19720 0 1 21493
box 0 0 1 1
use contact_30  contact_30_135
timestamp 1634918361
transform 1 0 19040 0 1 8709
box 0 0 1 1
use contact_30  contact_30_136
timestamp 1634918361
transform 1 0 19040 0 1 6941
box 0 0 1 1
use contact_30  contact_30_137
timestamp 1634918361
transform 1 0 15776 0 1 17957
box 0 0 1 1
use contact_30  contact_30_138
timestamp 1634918361
transform 1 0 15776 0 1 18501
box 0 0 1 1
use contact_30  contact_30_139
timestamp 1634918361
transform 1 0 14960 0 1 19997
box 0 0 1 1
use contact_30  contact_30_140
timestamp 1634918361
transform 1 0 14960 0 1 20269
box 0 0 1 1
use contact_30  contact_30_141
timestamp 1634918361
transform 1 0 14960 0 1 20405
box 0 0 1 1
use contact_30  contact_30_142
timestamp 1634918361
transform 1 0 14960 0 1 20677
box 0 0 1 1
use contact_30  contact_30_143
timestamp 1634918361
transform 1 0 15096 0 1 18365
box 0 0 1 1
use contact_30  contact_30_144
timestamp 1634918361
transform 1 0 15096 0 1 18637
box 0 0 1 1
use contact_30  contact_30_145
timestamp 1634918361
transform 1 0 14960 0 1 15237
box 0 0 1 1
use contact_30  contact_30_146
timestamp 1634918361
transform 1 0 14960 0 1 15509
box 0 0 1 1
use contact_30  contact_30_147
timestamp 1634918361
transform 1 0 15096 0 1 16325
box 0 0 1 1
use contact_30  contact_30_148
timestamp 1634918361
transform 1 0 15096 0 1 16053
box 0 0 1 1
use contact_30  contact_30_149
timestamp 1634918361
transform 1 0 14960 0 1 15645
box 0 0 1 1
use contact_30  contact_30_150
timestamp 1634918361
transform 1 0 14960 0 1 15917
box 0 0 1 1
use contact_30  contact_30_151
timestamp 1634918361
transform 1 0 15096 0 1 19861
box 0 0 1 1
use contact_30  contact_30_152
timestamp 1634918361
transform 1 0 15096 0 1 19589
box 0 0 1 1
use contact_30  contact_30_153
timestamp 1634918361
transform 1 0 15096 0 1 16461
box 0 0 1 1
use contact_30  contact_30_154
timestamp 1634918361
transform 1 0 15096 0 1 16733
box 0 0 1 1
use contact_30  contact_30_155
timestamp 1634918361
transform 1 0 15096 0 1 16869
box 0 0 1 1
use contact_30  contact_30_156
timestamp 1634918361
transform 1 0 15096 0 1 17141
box 0 0 1 1
use contact_30  contact_30_157
timestamp 1634918361
transform 1 0 14960 0 1 18773
box 0 0 1 1
use contact_30  contact_30_158
timestamp 1634918361
transform 1 0 14960 0 1 19045
box 0 0 1 1
use contact_30  contact_30_159
timestamp 1634918361
transform 1 0 14960 0 1 19453
box 0 0 1 1
use contact_30  contact_30_160
timestamp 1634918361
transform 1 0 14960 0 1 19181
box 0 0 1 1
use contact_30  contact_30_161
timestamp 1634918361
transform 1 0 14144 0 1 20405
box 0 0 1 1
use contact_30  contact_30_162
timestamp 1634918361
transform 1 0 14144 0 1 20677
box 0 0 1 1
use contact_30  contact_30_163
timestamp 1634918361
transform 1 0 14280 0 1 16053
box 0 0 1 1
use contact_30  contact_30_164
timestamp 1634918361
transform 1 0 14280 0 1 16325
box 0 0 1 1
use contact_30  contact_30_165
timestamp 1634918361
transform 1 0 14144 0 1 16733
box 0 0 1 1
use contact_30  contact_30_166
timestamp 1634918361
transform 1 0 14144 0 1 16461
box 0 0 1 1
use contact_30  contact_30_167
timestamp 1634918361
transform 1 0 14144 0 1 17549
box 0 0 1 1
use contact_30  contact_30_168
timestamp 1634918361
transform 1 0 14144 0 1 17277
box 0 0 1 1
use contact_30  contact_30_169
timestamp 1634918361
transform 1 0 14280 0 1 16869
box 0 0 1 1
use contact_30  contact_30_170
timestamp 1634918361
transform 1 0 14280 0 1 17141
box 0 0 1 1
use contact_30  contact_30_171
timestamp 1634918361
transform 1 0 14144 0 1 20269
box 0 0 1 1
use contact_30  contact_30_172
timestamp 1634918361
transform 1 0 14144 0 1 19997
box 0 0 1 1
use contact_30  contact_30_173
timestamp 1634918361
transform 1 0 14280 0 1 15917
box 0 0 1 1
use contact_30  contact_30_174
timestamp 1634918361
transform 1 0 14280 0 1 15645
box 0 0 1 1
use contact_30  contact_30_175
timestamp 1634918361
transform 1 0 14144 0 1 15237
box 0 0 1 1
use contact_30  contact_30_176
timestamp 1634918361
transform 1 0 14144 0 1 15509
box 0 0 1 1
use contact_30  contact_30_177
timestamp 1634918361
transform 1 0 14144 0 1 17685
box 0 0 1 1
use contact_30  contact_30_178
timestamp 1634918361
transform 1 0 14144 0 1 17957
box 0 0 1 1
use contact_30  contact_30_179
timestamp 1634918361
transform 1 0 14144 0 1 19181
box 0 0 1 1
use contact_30  contact_30_180
timestamp 1634918361
transform 1 0 14144 0 1 19453
box 0 0 1 1
use contact_30  contact_30_181
timestamp 1634918361
transform 1 0 14144 0 1 19861
box 0 0 1 1
use contact_30  contact_30_182
timestamp 1634918361
transform 1 0 14144 0 1 19589
box 0 0 1 1
use contact_30  contact_30_183
timestamp 1634918361
transform 1 0 12512 0 1 17685
box 0 0 1 1
use contact_30  contact_30_184
timestamp 1634918361
transform 1 0 12512 0 1 18229
box 0 0 1 1
use contact_30  contact_30_185
timestamp 1634918361
transform 1 0 12784 0 1 15645
box 0 0 1 1
use contact_30  contact_30_186
timestamp 1634918361
transform 1 0 12784 0 1 15917
box 0 0 1 1
use contact_30  contact_30_187
timestamp 1634918361
transform 1 0 12648 0 1 17413
box 0 0 1 1
use contact_30  contact_30_188
timestamp 1634918361
transform 1 0 12648 0 1 16053
box 0 0 1 1
use contact_30  contact_30_189
timestamp 1634918361
transform 1 0 12512 0 1 15101
box 0 0 1 1
use contact_30  contact_30_190
timestamp 1634918361
transform 1 0 12512 0 1 14829
box 0 0 1 1
use contact_30  contact_30_191
timestamp 1634918361
transform 1 0 12104 0 1 14829
box 0 0 1 1
use contact_30  contact_30_192
timestamp 1634918361
transform 1 0 12104 0 1 15101
box 0 0 1 1
use contact_30  contact_30_193
timestamp 1634918361
transform 1 0 11968 0 1 15917
box 0 0 1 1
use contact_30  contact_30_194
timestamp 1634918361
transform 1 0 11968 0 1 15237
box 0 0 1 1
use contact_30  contact_30_195
timestamp 1634918361
transform 1 0 11832 0 1 18229
box 0 0 1 1
use contact_30  contact_30_196
timestamp 1634918361
transform 1 0 11832 0 1 17685
box 0 0 1 1
use contact_30  contact_30_197
timestamp 1634918361
transform 1 0 9520 0 1 549
box 0 0 1 1
use contact_30  contact_30_198
timestamp 1634918361
transform 1 0 9520 0 1 2453
box 0 0 1 1
use contact_30  contact_30_199
timestamp 1634918361
transform 1 0 9248 0 1 2589
box 0 0 1 1
use contact_30  contact_30_200
timestamp 1634918361
transform 1 0 9248 0 1 5309
box 0 0 1 1
use contact_30  contact_30_201
timestamp 1634918361
transform 1 0 9520 0 1 8165
box 0 0 1 1
use contact_30  contact_30_202
timestamp 1634918361
transform 1 0 9384 0 1 5445
box 0 0 1 1
use contact_30  contact_30_203
timestamp 1634918361
transform 1 0 9520 0 1 8301
box 0 0 1 1
use contact_30  contact_30_204
timestamp 1634918361
transform 1 0 9520 0 1 11021
box 0 0 1 1
use contact_30  contact_30_205
timestamp 1634918361
transform 1 0 10472 0 1 15101
box 0 0 1 1
use contact_30  contact_30_206
timestamp 1634918361
transform 1 0 10472 0 1 14013
box 0 0 1 1
use contact_30  contact_30_207
timestamp 1634918361
transform 1 0 9520 0 1 11157
box 0 0 1 1
use contact_30  contact_30_208
timestamp 1634918361
transform 1 0 9520 0 1 13741
box 0 0 1 1
use contact_30  contact_30_209
timestamp 1634918361
transform 1 0 8840 0 1 26661
box 0 0 1 1
use contact_30  contact_30_210
timestamp 1634918361
transform 1 0 8840 0 1 24077
box 0 0 1 1
use contact_30  contact_30_211
timestamp 1634918361
transform 1 0 10472 0 1 17685
box 0 0 1 1
use contact_30  contact_30_212
timestamp 1634918361
transform 1 0 10472 0 1 21085
box 0 0 1 1
use contact_30  contact_30_213
timestamp 1634918361
transform 1 0 8840 0 1 23805
box 0 0 1 1
use contact_30  contact_30_214
timestamp 1634918361
transform 1 0 8840 0 1 21221
box 0 0 1 1
use contact_30  contact_30_215
timestamp 1634918361
transform 1 0 3944 0 1 20813
box 0 0 1 1
use contact_30  contact_30_216
timestamp 1634918361
transform 1 0 3944 0 1 18229
box 0 0 1 1
use contact_30  contact_30_217
timestamp 1634918361
transform 1 0 4080 0 1 9661
box 0 0 1 1
use contact_30  contact_30_218
timestamp 1634918361
transform 1 0 4080 0 1 12381
box 0 0 1 1
use contact_30  contact_30_219
timestamp 1634918361
transform 1 0 544 0 1 18093
box 0 0 1 1
use contact_30  contact_30_220
timestamp 1634918361
transform 1 0 3808 0 1 15373
box 0 0 1 1
use contact_30  contact_30_221
timestamp 1634918361
transform 1 0 3808 0 1 18093
box 0 0 1 1
use contact_30  contact_30_222
timestamp 1634918361
transform 1 0 3400 0 1 12517
box 0 0 1 1
use contact_30  contact_30_223
timestamp 1634918361
transform 1 0 3400 0 1 15237
box 0 0 1 1
use contact_30  contact_30_224
timestamp 1634918361
transform 1 0 544 0 1 5581
box 0 0 1 1
use contact_30  contact_30_225
timestamp 1634918361
transform 1 0 544 0 1 2453
box 0 0 1 1
use contact_30  contact_30_226
timestamp 1634918361
transform 1 0 42160 0 1 3813
box 0 0 1 1
use contact_30  contact_30_227
timestamp 1634918361
transform 1 0 42160 0 1 22173
box 0 0 1 1
use contact_30  contact_30_228
timestamp 1634918361
transform 1 0 42160 0 1 17141
box 0 0 1 1
use contact_30  contact_30_229
timestamp 1634918361
transform 1 0 42160 0 1 30741
box 0 0 1 1
use contact_30  contact_30_230
timestamp 1634918361
transform 1 0 42160 0 1 8709
box 0 0 1 1
use contact_30  contact_30_231
timestamp 1634918361
transform 1 0 42160 0 1 2045
box 0 0 1 1
use contact_30  contact_30_232
timestamp 1634918361
transform 1 0 42160 0 1 28837
box 0 0 1 1
use contact_30  contact_30_233
timestamp 1634918361
transform 1 0 42160 0 1 12245
box 0 0 1 1
use contact_30  contact_30_234
timestamp 1634918361
transform 1 0 42160 0 1 27341
box 0 0 1 1
use contact_30  contact_30_235
timestamp 1634918361
transform 1 0 42160 0 1 18909
box 0 0 1 1
use contact_30  contact_30_236
timestamp 1634918361
transform 1 0 42160 0 1 23805
box 0 0 1 1
use contact_30  contact_30_237
timestamp 1634918361
transform 1 0 42160 0 1 10341
box 0 0 1 1
use contact_30  contact_30_238
timestamp 1634918361
transform 1 0 42160 0 1 13741
box 0 0 1 1
use contact_30  contact_30_239
timestamp 1634918361
transform 1 0 42160 0 1 15373
box 0 0 1 1
use contact_30  contact_30_240
timestamp 1634918361
transform 1 0 42160 0 1 7077
box 0 0 1 1
use contact_30  contact_30_241
timestamp 1634918361
transform 1 0 42160 0 1 5309
box 0 0 1 1
use contact_30  contact_30_242
timestamp 1634918361
transform 1 0 42160 0 1 20405
box 0 0 1 1
use contact_30  contact_30_243
timestamp 1634918361
transform 1 0 42160 0 1 25437
box 0 0 1 1
use contact_30  contact_30_244
timestamp 1634918361
transform 1 0 40664 0 1 31829
box 0 0 1 1
use contact_30  contact_30_245
timestamp 1634918361
transform 1 0 40664 0 1 31421
box 0 0 1 1
use contact_30  contact_30_246
timestamp 1634918361
transform 1 0 40800 0 1 1229
box 0 0 1 1
use contact_30  contact_30_247
timestamp 1634918361
transform 1 0 40800 0 1 1637
box 0 0 1 1
use contact_30  contact_30_248
timestamp 1634918361
transform 1 0 41616 0 1 18909
box 0 0 1 1
use contact_30  contact_30_249
timestamp 1634918361
transform 1 0 41616 0 1 19181
box 0 0 1 1
use contact_30  contact_30_250
timestamp 1634918361
transform 1 0 41616 0 1 17141
box 0 0 1 1
use contact_30  contact_30_251
timestamp 1634918361
transform 1 0 41616 0 1 16461
box 0 0 1 1
use contact_30  contact_30_252
timestamp 1634918361
transform 1 0 41616 0 1 23941
box 0 0 1 1
use contact_30  contact_30_253
timestamp 1634918361
transform 1 0 41616 0 1 24757
box 0 0 1 1
use contact_30  contact_30_254
timestamp 1634918361
transform 1 0 39032 0 1 1229
box 0 0 1 1
use contact_30  contact_30_255
timestamp 1634918361
transform 1 0 39032 0 1 1637
box 0 0 1 1
use contact_30  contact_30_256
timestamp 1634918361
transform 1 0 38896 0 1 31829
box 0 0 1 1
use contact_30  contact_30_257
timestamp 1634918361
transform 1 0 38896 0 1 31421
box 0 0 1 1
use contact_30  contact_30_258
timestamp 1634918361
transform 1 0 37400 0 1 1229
box 0 0 1 1
use contact_30  contact_30_259
timestamp 1634918361
transform 1 0 37400 0 1 1637
box 0 0 1 1
use contact_30  contact_30_260
timestamp 1634918361
transform 1 0 37264 0 1 31829
box 0 0 1 1
use contact_30  contact_30_261
timestamp 1634918361
transform 1 0 37264 0 1 31421
box 0 0 1 1
use contact_30  contact_30_262
timestamp 1634918361
transform 1 0 35632 0 1 31829
box 0 0 1 1
use contact_30  contact_30_263
timestamp 1634918361
transform 1 0 35632 0 1 31421
box 0 0 1 1
use contact_30  contact_30_264
timestamp 1634918361
transform 1 0 35632 0 1 1229
box 0 0 1 1
use contact_30  contact_30_265
timestamp 1634918361
transform 1 0 35632 0 1 1637
box 0 0 1 1
use contact_30  contact_30_266
timestamp 1634918361
transform 1 0 34816 0 1 13333
box 0 0 1 1
use contact_30  contact_30_267
timestamp 1634918361
transform 1 0 34816 0 1 10613
box 0 0 1 1
use contact_30  contact_30_268
timestamp 1634918361
transform 1 0 34272 0 1 28973
box 0 0 1 1
use contact_30  contact_30_269
timestamp 1634918361
transform 1 0 34272 0 1 26389
box 0 0 1 1
use contact_30  contact_30_270
timestamp 1634918361
transform 1 0 34136 0 1 26253
box 0 0 1 1
use contact_30  contact_30_271
timestamp 1634918361
transform 1 0 34136 0 1 23533
box 0 0 1 1
use contact_30  contact_30_272
timestamp 1634918361
transform 1 0 34000 0 1 31829
box 0 0 1 1
use contact_30  contact_30_273
timestamp 1634918361
transform 1 0 34000 0 1 31421
box 0 0 1 1
use contact_30  contact_30_274
timestamp 1634918361
transform 1 0 34136 0 1 29109
box 0 0 1 1
use contact_30  contact_30_275
timestamp 1634918361
transform 1 0 34136 0 1 31285
box 0 0 1 1
use contact_30  contact_30_276
timestamp 1634918361
transform 1 0 34000 0 1 1229
box 0 0 1 1
use contact_30  contact_30_277
timestamp 1634918361
transform 1 0 34000 0 1 1637
box 0 0 1 1
use contact_30  contact_30_278
timestamp 1634918361
transform 1 0 32776 0 1 13469
box 0 0 1 1
use contact_30  contact_30_279
timestamp 1634918361
transform 1 0 32776 0 1 15101
box 0 0 1 1
use contact_30  contact_30_280
timestamp 1634918361
transform 1 0 32232 0 1 1229
box 0 0 1 1
use contact_30  contact_30_281
timestamp 1634918361
transform 1 0 32232 0 1 1637
box 0 0 1 1
use contact_30  contact_30_282
timestamp 1634918361
transform 1 0 32232 0 1 31829
box 0 0 1 1
use contact_30  contact_30_283
timestamp 1634918361
transform 1 0 32232 0 1 31421
box 0 0 1 1
use contact_30  contact_30_284
timestamp 1634918361
transform 1 0 31280 0 1 15917
box 0 0 1 1
use contact_30  contact_30_285
timestamp 1634918361
transform 1 0 31280 0 1 15237
box 0 0 1 1
use contact_30  contact_30_286
timestamp 1634918361
transform 1 0 31144 0 1 17685
box 0 0 1 1
use contact_30  contact_30_287
timestamp 1634918361
transform 1 0 31144 0 1 18229
box 0 0 1 1
use contact_30  contact_30_288
timestamp 1634918361
transform 1 0 30600 0 1 31829
box 0 0 1 1
use contact_30  contact_30_289
timestamp 1634918361
transform 1 0 30600 0 1 31421
box 0 0 1 1
use contact_30  contact_30_290
timestamp 1634918361
transform 1 0 30600 0 1 1229
box 0 0 1 1
use contact_30  contact_30_291
timestamp 1634918361
transform 1 0 30600 0 1 1637
box 0 0 1 1
use contact_30  contact_30_292
timestamp 1634918361
transform 1 0 30464 0 1 16053
box 0 0 1 1
use contact_30  contact_30_293
timestamp 1634918361
transform 1 0 30464 0 1 17413
box 0 0 1 1
use contact_30  contact_30_294
timestamp 1634918361
transform 1 0 30464 0 1 17685
box 0 0 1 1
use contact_30  contact_30_295
timestamp 1634918361
transform 1 0 30464 0 1 18229
box 0 0 1 1
use contact_30  contact_30_296
timestamp 1634918361
transform 1 0 28968 0 1 31829
box 0 0 1 1
use contact_30  contact_30_297
timestamp 1634918361
transform 1 0 28968 0 1 31421
box 0 0 1 1
use contact_30  contact_30_298
timestamp 1634918361
transform 1 0 28968 0 1 1229
box 0 0 1 1
use contact_30  contact_30_299
timestamp 1634918361
transform 1 0 28968 0 1 1637
box 0 0 1 1
use contact_30  contact_30_300
timestamp 1634918361
transform 1 0 28968 0 1 16461
box 0 0 1 1
use contact_30  contact_30_301
timestamp 1634918361
transform 1 0 28968 0 1 16733
box 0 0 1 1
use contact_30  contact_30_302
timestamp 1634918361
transform 1 0 28968 0 1 16869
box 0 0 1 1
use contact_30  contact_30_303
timestamp 1634918361
transform 1 0 28968 0 1 17141
box 0 0 1 1
use contact_30  contact_30_304
timestamp 1634918361
transform 1 0 28968 0 1 15509
box 0 0 1 1
use contact_30  contact_30_305
timestamp 1634918361
transform 1 0 28968 0 1 15237
box 0 0 1 1
use contact_30  contact_30_306
timestamp 1634918361
transform 1 0 28968 0 1 17277
box 0 0 1 1
use contact_30  contact_30_307
timestamp 1634918361
transform 1 0 28968 0 1 17549
box 0 0 1 1
use contact_30  contact_30_308
timestamp 1634918361
transform 1 0 28968 0 1 20677
box 0 0 1 1
use contact_30  contact_30_309
timestamp 1634918361
transform 1 0 28968 0 1 20405
box 0 0 1 1
use contact_30  contact_30_310
timestamp 1634918361
transform 1 0 28968 0 1 15645
box 0 0 1 1
use contact_30  contact_30_311
timestamp 1634918361
transform 1 0 28968 0 1 15917
box 0 0 1 1
use contact_30  contact_30_312
timestamp 1634918361
transform 1 0 28968 0 1 16325
box 0 0 1 1
use contact_30  contact_30_313
timestamp 1634918361
transform 1 0 28968 0 1 16053
box 0 0 1 1
use contact_30  contact_30_314
timestamp 1634918361
transform 1 0 28832 0 1 19589
box 0 0 1 1
use contact_30  contact_30_315
timestamp 1634918361
transform 1 0 28832 0 1 19861
box 0 0 1 1
use contact_30  contact_30_316
timestamp 1634918361
transform 1 0 28968 0 1 20269
box 0 0 1 1
use contact_30  contact_30_317
timestamp 1634918361
transform 1 0 28968 0 1 19997
box 0 0 1 1
use contact_30  contact_30_318
timestamp 1634918361
transform 1 0 28968 0 1 17685
box 0 0 1 1
use contact_30  contact_30_319
timestamp 1634918361
transform 1 0 28968 0 1 17957
box 0 0 1 1
use contact_30  contact_30_320
timestamp 1634918361
transform 1 0 28832 0 1 19453
box 0 0 1 1
use contact_30  contact_30_321
timestamp 1634918361
transform 1 0 28832 0 1 19181
box 0 0 1 1
use contact_30  contact_30_322
timestamp 1634918361
transform 1 0 28016 0 1 19045
box 0 0 1 1
use contact_30  contact_30_323
timestamp 1634918361
transform 1 0 28016 0 1 18773
box 0 0 1 1
use contact_30  contact_30_324
timestamp 1634918361
transform 1 0 28016 0 1 20405
box 0 0 1 1
use contact_30  contact_30_325
timestamp 1634918361
transform 1 0 28016 0 1 20677
box 0 0 1 1
use contact_30  contact_30_326
timestamp 1634918361
transform 1 0 28152 0 1 15645
box 0 0 1 1
use contact_30  contact_30_327
timestamp 1634918361
transform 1 0 28152 0 1 15917
box 0 0 1 1
use contact_30  contact_30_328
timestamp 1634918361
transform 1 0 28152 0 1 18637
box 0 0 1 1
use contact_30  contact_30_329
timestamp 1634918361
transform 1 0 28152 0 1 18365
box 0 0 1 1
use contact_30  contact_30_330
timestamp 1634918361
transform 1 0 28288 0 1 16053
box 0 0 1 1
use contact_30  contact_30_331
timestamp 1634918361
transform 1 0 28288 0 1 16325
box 0 0 1 1
use contact_30  contact_30_332
timestamp 1634918361
transform 1 0 28152 0 1 19181
box 0 0 1 1
use contact_30  contact_30_333
timestamp 1634918361
transform 1 0 28152 0 1 19453
box 0 0 1 1
use contact_30  contact_30_334
timestamp 1634918361
transform 1 0 28152 0 1 17141
box 0 0 1 1
use contact_30  contact_30_335
timestamp 1634918361
transform 1 0 28152 0 1 16869
box 0 0 1 1
use contact_30  contact_30_336
timestamp 1634918361
transform 1 0 28152 0 1 16461
box 0 0 1 1
use contact_30  contact_30_337
timestamp 1634918361
transform 1 0 28152 0 1 16733
box 0 0 1 1
use contact_30  contact_30_338
timestamp 1634918361
transform 1 0 28016 0 1 20269
box 0 0 1 1
use contact_30  contact_30_339
timestamp 1634918361
transform 1 0 28016 0 1 19997
box 0 0 1 1
use contact_30  contact_30_340
timestamp 1634918361
transform 1 0 28288 0 1 19589
box 0 0 1 1
use contact_30  contact_30_341
timestamp 1634918361
transform 1 0 28288 0 1 19861
box 0 0 1 1
use contact_30  contact_30_342
timestamp 1634918361
transform 1 0 28016 0 1 15509
box 0 0 1 1
use contact_30  contact_30_343
timestamp 1634918361
transform 1 0 28016 0 1 15237
box 0 0 1 1
use contact_30  contact_30_344
timestamp 1634918361
transform 1 0 28016 0 1 20813
box 0 0 1 1
use contact_30  contact_30_345
timestamp 1634918361
transform 1 0 28016 0 1 21221
box 0 0 1 1
use contact_30  contact_30_346
timestamp 1634918361
transform 1 0 27880 0 1 20813
box 0 0 1 1
use contact_30  contact_30_347
timestamp 1634918361
transform 1 0 27880 0 1 21221
box 0 0 1 1
use contact_30  contact_30_348
timestamp 1634918361
transform 1 0 27200 0 1 31829
box 0 0 1 1
use contact_30  contact_30_349
timestamp 1634918361
transform 1 0 27200 0 1 31421
box 0 0 1 1
use contact_30  contact_30_350
timestamp 1634918361
transform 1 0 27336 0 1 1229
box 0 0 1 1
use contact_30  contact_30_351
timestamp 1634918361
transform 1 0 27336 0 1 1637
box 0 0 1 1
use contact_30  contact_30_352
timestamp 1634918361
transform 1 0 25432 0 1 1229
box 0 0 1 1
use contact_30  contact_30_353
timestamp 1634918361
transform 1 0 25432 0 1 1637
box 0 0 1 1
use contact_30  contact_30_354
timestamp 1634918361
transform 1 0 25568 0 1 31829
box 0 0 1 1
use contact_30  contact_30_355
timestamp 1634918361
transform 1 0 25568 0 1 31421
box 0 0 1 1
use contact_30  contact_30_356
timestamp 1634918361
transform 1 0 26248 0 1 21357
box 0 0 1 1
use contact_30  contact_30_357
timestamp 1634918361
transform 1 0 26248 0 1 21629
box 0 0 1 1
use contact_30  contact_30_358
timestamp 1634918361
transform 1 0 24344 0 1 22173
box 0 0 1 1
use contact_30  contact_30_359
timestamp 1634918361
transform 1 0 24344 0 1 21765
box 0 0 1 1
use contact_30  contact_30_360
timestamp 1634918361
transform 1 0 24072 0 1 22173
box 0 0 1 1
use contact_30  contact_30_361
timestamp 1634918361
transform 1 0 24072 0 1 21765
box 0 0 1 1
use contact_30  contact_30_362
timestamp 1634918361
transform 1 0 23936 0 1 13741
box 0 0 1 1
use contact_30  contact_30_363
timestamp 1634918361
transform 1 0 23936 0 1 14149
box 0 0 1 1
use contact_30  contact_30_364
timestamp 1634918361
transform 1 0 23800 0 1 31829
box 0 0 1 1
use contact_30  contact_30_365
timestamp 1634918361
transform 1 0 23800 0 1 31421
box 0 0 1 1
use contact_30  contact_30_366
timestamp 1634918361
transform 1 0 23528 0 1 1229
box 0 0 1 1
use contact_30  contact_30_367
timestamp 1634918361
transform 1 0 23528 0 1 1637
box 0 0 1 1
use contact_30  contact_30_368
timestamp 1634918361
transform 1 0 24344 0 1 8029
box 0 0 1 1
use contact_30  contact_30_369
timestamp 1634918361
transform 1 0 24344 0 1 8437
box 0 0 1 1
use contact_30  contact_30_370
timestamp 1634918361
transform 1 0 23800 0 1 13741
box 0 0 1 1
use contact_30  contact_30_371
timestamp 1634918361
transform 1 0 23800 0 1 14149
box 0 0 1 1
use contact_30  contact_30_372
timestamp 1634918361
transform 1 0 23256 0 1 14149
box 0 0 1 1
use contact_30  contact_30_373
timestamp 1634918361
transform 1 0 23256 0 1 13741
box 0 0 1 1
use contact_30  contact_30_374
timestamp 1634918361
transform 1 0 23256 0 1 21765
box 0 0 1 1
use contact_30  contact_30_375
timestamp 1634918361
transform 1 0 23256 0 1 22173
box 0 0 1 1
use contact_30  contact_30_376
timestamp 1634918361
transform 1 0 23120 0 1 13741
box 0 0 1 1
use contact_30  contact_30_377
timestamp 1634918361
transform 1 0 23120 0 1 14149
box 0 0 1 1
use contact_30  contact_30_378
timestamp 1634918361
transform 1 0 22712 0 1 13741
box 0 0 1 1
use contact_30  contact_30_379
timestamp 1634918361
transform 1 0 22712 0 1 14149
box 0 0 1 1
use contact_30  contact_30_380
timestamp 1634918361
transform 1 0 22712 0 1 22173
box 0 0 1 1
use contact_30  contact_30_381
timestamp 1634918361
transform 1 0 22712 0 1 21765
box 0 0 1 1
use contact_30  contact_30_382
timestamp 1634918361
transform 1 0 22576 0 1 24213
box 0 0 1 1
use contact_30  contact_30_383
timestamp 1634918361
transform 1 0 22576 0 1 24893
box 0 0 1 1
use contact_30  contact_30_384
timestamp 1634918361
transform 1 0 22304 0 1 31829
box 0 0 1 1
use contact_30  contact_30_385
timestamp 1634918361
transform 1 0 22304 0 1 31421
box 0 0 1 1
use contact_30  contact_30_386
timestamp 1634918361
transform 1 0 22304 0 1 1229
box 0 0 1 1
use contact_30  contact_30_387
timestamp 1634918361
transform 1 0 22304 0 1 1637
box 0 0 1 1
use contact_30  contact_30_388
timestamp 1634918361
transform 1 0 22576 0 1 11837
box 0 0 1 1
use contact_30  contact_30_389
timestamp 1634918361
transform 1 0 22576 0 1 13605
box 0 0 1 1
use contact_30  contact_30_390
timestamp 1634918361
transform 1 0 22032 0 1 14149
box 0 0 1 1
use contact_30  contact_30_391
timestamp 1634918361
transform 1 0 22032 0 1 13741
box 0 0 1 1
use contact_30  contact_30_392
timestamp 1634918361
transform 1 0 22032 0 1 21765
box 0 0 1 1
use contact_30  contact_30_393
timestamp 1634918361
transform 1 0 22032 0 1 22173
box 0 0 1 1
use contact_30  contact_30_394
timestamp 1634918361
transform 1 0 21488 0 1 13741
box 0 0 1 1
use contact_30  contact_30_395
timestamp 1634918361
transform 1 0 21488 0 1 14149
box 0 0 1 1
use contact_30  contact_30_396
timestamp 1634918361
transform 1 0 21488 0 1 24213
box 0 0 1 1
use contact_30  contact_30_397
timestamp 1634918361
transform 1 0 21488 0 1 24893
box 0 0 1 1
use contact_30  contact_30_398
timestamp 1634918361
transform 1 0 20672 0 1 8437
box 0 0 1 1
use contact_30  contact_30_399
timestamp 1634918361
transform 1 0 20672 0 1 9253
box 0 0 1 1
use contact_30  contact_30_400
timestamp 1634918361
transform 1 0 20808 0 1 14149
box 0 0 1 1
use contact_30  contact_30_401
timestamp 1634918361
transform 1 0 20808 0 1 13741
box 0 0 1 1
use contact_30  contact_30_402
timestamp 1634918361
transform 1 0 20808 0 1 21765
box 0 0 1 1
use contact_30  contact_30_403
timestamp 1634918361
transform 1 0 20808 0 1 22173
box 0 0 1 1
use contact_30  contact_30_404
timestamp 1634918361
transform 1 0 20672 0 1 1229
box 0 0 1 1
use contact_30  contact_30_405
timestamp 1634918361
transform 1 0 20672 0 1 1637
box 0 0 1 1
use contact_30  contact_30_406
timestamp 1634918361
transform 1 0 20264 0 1 31829
box 0 0 1 1
use contact_30  contact_30_407
timestamp 1634918361
transform 1 0 20264 0 1 31421
box 0 0 1 1
use contact_30  contact_30_408
timestamp 1634918361
transform 1 0 20264 0 1 22173
box 0 0 1 1
use contact_30  contact_30_409
timestamp 1634918361
transform 1 0 20264 0 1 21765
box 0 0 1 1
use contact_30  contact_30_410
timestamp 1634918361
transform 1 0 20264 0 1 11701
box 0 0 1 1
use contact_30  contact_30_411
timestamp 1634918361
transform 1 0 20264 0 1 11021
box 0 0 1 1
use contact_30  contact_30_412
timestamp 1634918361
transform 1 0 19992 0 1 10885
box 0 0 1 1
use contact_30  contact_30_413
timestamp 1634918361
transform 1 0 19992 0 1 9525
box 0 0 1 1
use contact_30  contact_30_414
timestamp 1634918361
transform 1 0 19584 0 1 24077
box 0 0 1 1
use contact_30  contact_30_415
timestamp 1634918361
transform 1 0 19584 0 1 22309
box 0 0 1 1
use contact_30  contact_30_416
timestamp 1634918361
transform 1 0 19584 0 1 21765
box 0 0 1 1
use contact_30  contact_30_417
timestamp 1634918361
transform 1 0 19584 0 1 22173
box 0 0 1 1
use contact_30  contact_30_418
timestamp 1634918361
transform 1 0 19040 0 1 13741
box 0 0 1 1
use contact_30  contact_30_419
timestamp 1634918361
transform 1 0 19040 0 1 14149
box 0 0 1 1
use contact_30  contact_30_420
timestamp 1634918361
transform 1 0 18768 0 1 1229
box 0 0 1 1
use contact_30  contact_30_421
timestamp 1634918361
transform 1 0 18768 0 1 1637
box 0 0 1 1
use contact_30  contact_30_422
timestamp 1634918361
transform 1 0 18768 0 1 31829
box 0 0 1 1
use contact_30  contact_30_423
timestamp 1634918361
transform 1 0 18768 0 1 31421
box 0 0 1 1
use contact_30  contact_30_424
timestamp 1634918361
transform 1 0 19312 0 1 8437
box 0 0 1 1
use contact_30  contact_30_425
timestamp 1634918361
transform 1 0 19312 0 1 8029
box 0 0 1 1
use contact_30  contact_30_426
timestamp 1634918361
transform 1 0 17680 0 1 14285
box 0 0 1 1
use contact_30  contact_30_427
timestamp 1634918361
transform 1 0 17680 0 1 14557
box 0 0 1 1
use contact_30  contact_30_428
timestamp 1634918361
transform 1 0 17272 0 1 1229
box 0 0 1 1
use contact_30  contact_30_429
timestamp 1634918361
transform 1 0 17272 0 1 1637
box 0 0 1 1
use contact_30  contact_30_430
timestamp 1634918361
transform 1 0 17272 0 1 31829
box 0 0 1 1
use contact_30  contact_30_431
timestamp 1634918361
transform 1 0 17272 0 1 31421
box 0 0 1 1
use contact_30  contact_30_432
timestamp 1634918361
transform 1 0 15368 0 1 1229
box 0 0 1 1
use contact_30  contact_30_433
timestamp 1634918361
transform 1 0 15368 0 1 1637
box 0 0 1 1
use contact_30  contact_30_434
timestamp 1634918361
transform 1 0 15640 0 1 31829
box 0 0 1 1
use contact_30  contact_30_435
timestamp 1634918361
transform 1 0 15640 0 1 31421
box 0 0 1 1
use contact_30  contact_30_436
timestamp 1634918361
transform 1 0 15232 0 1 19453
box 0 0 1 1
use contact_30  contact_30_437
timestamp 1634918361
transform 1 0 15232 0 1 19181
box 0 0 1 1
use contact_30  contact_30_438
timestamp 1634918361
transform 1 0 15232 0 1 17141
box 0 0 1 1
use contact_30  contact_30_439
timestamp 1634918361
transform 1 0 15232 0 1 16869
box 0 0 1 1
use contact_30  contact_30_440
timestamp 1634918361
transform 1 0 18088 0 1 21629
box 0 0 1 1
use contact_30  contact_30_441
timestamp 1634918361
transform 1 0 18088 0 1 20813
box 0 0 1 1
use contact_30  contact_30_442
timestamp 1634918361
transform 1 0 16184 0 1 17957
box 0 0 1 1
use contact_30  contact_30_443
timestamp 1634918361
transform 1 0 16184 0 1 18229
box 0 0 1 1
use contact_30  contact_30_444
timestamp 1634918361
transform 1 0 15232 0 1 19045
box 0 0 1 1
use contact_30  contact_30_445
timestamp 1634918361
transform 1 0 15232 0 1 18773
box 0 0 1 1
use contact_30  contact_30_446
timestamp 1634918361
transform 1 0 15368 0 1 18365
box 0 0 1 1
use contact_30  contact_30_447
timestamp 1634918361
transform 1 0 15368 0 1 18637
box 0 0 1 1
use contact_30  contact_30_448
timestamp 1634918361
transform 1 0 15232 0 1 19589
box 0 0 1 1
use contact_30  contact_30_449
timestamp 1634918361
transform 1 0 15232 0 1 19861
box 0 0 1 1
use contact_30  contact_30_450
timestamp 1634918361
transform 1 0 15368 0 1 14693
box 0 0 1 1
use contact_30  contact_30_451
timestamp 1634918361
transform 1 0 15368 0 1 15101
box 0 0 1 1
use contact_30  contact_30_452
timestamp 1634918361
transform 1 0 15504 0 1 16733
box 0 0 1 1
use contact_30  contact_30_453
timestamp 1634918361
transform 1 0 15504 0 1 16461
box 0 0 1 1
use contact_30  contact_30_454
timestamp 1634918361
transform 1 0 15504 0 1 16053
box 0 0 1 1
use contact_30  contact_30_455
timestamp 1634918361
transform 1 0 15504 0 1 16325
box 0 0 1 1
use contact_30  contact_30_456
timestamp 1634918361
transform 1 0 15504 0 1 15917
box 0 0 1 1
use contact_30  contact_30_457
timestamp 1634918361
transform 1 0 15504 0 1 15645
box 0 0 1 1
use contact_30  contact_30_458
timestamp 1634918361
transform 1 0 15232 0 1 15237
box 0 0 1 1
use contact_30  contact_30_459
timestamp 1634918361
transform 1 0 15232 0 1 15509
box 0 0 1 1
use contact_30  contact_30_460
timestamp 1634918361
transform 1 0 15232 0 1 20677
box 0 0 1 1
use contact_30  contact_30_461
timestamp 1634918361
transform 1 0 15232 0 1 20405
box 0 0 1 1
use contact_30  contact_30_462
timestamp 1634918361
transform 1 0 15232 0 1 19997
box 0 0 1 1
use contact_30  contact_30_463
timestamp 1634918361
transform 1 0 15232 0 1 20269
box 0 0 1 1
use contact_30  contact_30_464
timestamp 1634918361
transform 1 0 14688 0 1 20677
box 0 0 1 1
use contact_30  contact_30_465
timestamp 1634918361
transform 1 0 14688 0 1 20405
box 0 0 1 1
use contact_30  contact_30_466
timestamp 1634918361
transform 1 0 14688 0 1 20269
box 0 0 1 1
use contact_30  contact_30_467
timestamp 1634918361
transform 1 0 14688 0 1 19997
box 0 0 1 1
use contact_30  contact_30_468
timestamp 1634918361
transform 1 0 14552 0 1 19589
box 0 0 1 1
use contact_30  contact_30_469
timestamp 1634918361
transform 1 0 14552 0 1 19861
box 0 0 1 1
use contact_30  contact_30_470
timestamp 1634918361
transform 1 0 14688 0 1 15509
box 0 0 1 1
use contact_30  contact_30_471
timestamp 1634918361
transform 1 0 14688 0 1 15237
box 0 0 1 1
use contact_30  contact_30_472
timestamp 1634918361
transform 1 0 14552 0 1 19453
box 0 0 1 1
use contact_30  contact_30_473
timestamp 1634918361
transform 1 0 14552 0 1 19181
box 0 0 1 1
use contact_30  contact_30_474
timestamp 1634918361
transform 1 0 14552 0 1 16461
box 0 0 1 1
use contact_30  contact_30_475
timestamp 1634918361
transform 1 0 14552 0 1 16733
box 0 0 1 1
use contact_30  contact_30_476
timestamp 1634918361
transform 1 0 14688 0 1 17141
box 0 0 1 1
use contact_30  contact_30_477
timestamp 1634918361
transform 1 0 14688 0 1 16869
box 0 0 1 1
use contact_30  contact_30_478
timestamp 1634918361
transform 1 0 14688 0 1 16325
box 0 0 1 1
use contact_30  contact_30_479
timestamp 1634918361
transform 1 0 14688 0 1 16053
box 0 0 1 1
use contact_30  contact_30_480
timestamp 1634918361
transform 1 0 14688 0 1 15645
box 0 0 1 1
use contact_30  contact_30_481
timestamp 1634918361
transform 1 0 14688 0 1 15917
box 0 0 1 1
use contact_30  contact_30_482
timestamp 1634918361
transform 1 0 14688 0 1 17277
box 0 0 1 1
use contact_30  contact_30_483
timestamp 1634918361
transform 1 0 14688 0 1 17549
box 0 0 1 1
use contact_30  contact_30_484
timestamp 1634918361
transform 1 0 14688 0 1 17957
box 0 0 1 1
use contact_30  contact_30_485
timestamp 1634918361
transform 1 0 14688 0 1 17685
box 0 0 1 1
use contact_30  contact_30_486
timestamp 1634918361
transform 1 0 13736 0 1 1229
box 0 0 1 1
use contact_30  contact_30_487
timestamp 1634918361
transform 1 0 13736 0 1 1637
box 0 0 1 1
use contact_30  contact_30_488
timestamp 1634918361
transform 1 0 13736 0 1 31829
box 0 0 1 1
use contact_30  contact_30_489
timestamp 1634918361
transform 1 0 13736 0 1 31421
box 0 0 1 1
use contact_30  contact_30_490
timestamp 1634918361
transform 1 0 13056 0 1 17413
box 0 0 1 1
use contact_30  contact_30_491
timestamp 1634918361
transform 1 0 13056 0 1 16053
box 0 0 1 1
use contact_30  contact_30_492
timestamp 1634918361
transform 1 0 12376 0 1 17685
box 0 0 1 1
use contact_30  contact_30_493
timestamp 1634918361
transform 1 0 12376 0 1 18229
box 0 0 1 1
use contact_30  contact_30_494
timestamp 1634918361
transform 1 0 12240 0 1 15917
box 0 0 1 1
use contact_30  contact_30_495
timestamp 1634918361
transform 1 0 12240 0 1 15237
box 0 0 1 1
use contact_30  contact_30_496
timestamp 1634918361
transform 1 0 12104 0 1 31829
box 0 0 1 1
use contact_30  contact_30_497
timestamp 1634918361
transform 1 0 12104 0 1 31421
box 0 0 1 1
use contact_30  contact_30_498
timestamp 1634918361
transform 1 0 12240 0 1 1229
box 0 0 1 1
use contact_30  contact_30_499
timestamp 1634918361
transform 1 0 12240 0 1 1637
box 0 0 1 1
use contact_30  contact_30_500
timestamp 1634918361
transform 1 0 12240 0 1 18229
box 0 0 1 1
use contact_30  contact_30_501
timestamp 1634918361
transform 1 0 12240 0 1 17413
box 0 0 1 1
use contact_30  contact_30_502
timestamp 1634918361
transform 1 0 10336 0 1 1229
box 0 0 1 1
use contact_30  contact_30_503
timestamp 1634918361
transform 1 0 10336 0 1 1637
box 0 0 1 1
use contact_30  contact_30_504
timestamp 1634918361
transform 1 0 10336 0 1 31829
box 0 0 1 1
use contact_30  contact_30_505
timestamp 1634918361
transform 1 0 10336 0 1 31421
box 0 0 1 1
use contact_30  contact_30_506
timestamp 1634918361
transform 1 0 10880 0 1 15101
box 0 0 1 1
use contact_30  contact_30_507
timestamp 1634918361
transform 1 0 10880 0 1 12517
box 0 0 1 1
use contact_30  contact_30_508
timestamp 1634918361
transform 1 0 9384 0 1 12381
box 0 0 1 1
use contact_30  contact_30_509
timestamp 1634918361
transform 1 0 9384 0 1 9661
box 0 0 1 1
use contact_30  contact_30_510
timestamp 1634918361
transform 1 0 9520 0 1 4085
box 0 0 1 1
use contact_30  contact_30_511
timestamp 1634918361
transform 1 0 9520 0 1 6669
box 0 0 1 1
use contact_30  contact_30_512
timestamp 1634918361
transform 1 0 9384 0 1 9525
box 0 0 1 1
use contact_30  contact_30_513
timestamp 1634918361
transform 1 0 9384 0 1 6941
box 0 0 1 1
use contact_30  contact_30_514
timestamp 1634918361
transform 1 0 12240 0 1 18501
box 0 0 1 1
use contact_30  contact_30_515
timestamp 1634918361
transform 1 0 12240 0 1 22445
box 0 0 1 1
use contact_30  contact_30_516
timestamp 1634918361
transform 1 0 8976 0 1 25301
box 0 0 1 1
use contact_30  contact_30_517
timestamp 1634918361
transform 1 0 8976 0 1 22581
box 0 0 1 1
use contact_30  contact_30_518
timestamp 1634918361
transform 1 0 8704 0 1 1229
box 0 0 1 1
use contact_30  contact_30_519
timestamp 1634918361
transform 1 0 8704 0 1 1637
box 0 0 1 1
use contact_30  contact_30_520
timestamp 1634918361
transform 1 0 9384 0 1 3949
box 0 0 1 1
use contact_30  contact_30_521
timestamp 1634918361
transform 1 0 9384 0 1 1773
box 0 0 1 1
use contact_30  contact_30_522
timestamp 1634918361
transform 1 0 8704 0 1 31829
box 0 0 1 1
use contact_30  contact_30_523
timestamp 1634918361
transform 1 0 8704 0 1 31421
box 0 0 1 1
use contact_30  contact_30_524
timestamp 1634918361
transform 1 0 7072 0 1 31829
box 0 0 1 1
use contact_30  contact_30_525
timestamp 1634918361
transform 1 0 7072 0 1 31421
box 0 0 1 1
use contact_30  contact_30_526
timestamp 1634918361
transform 1 0 7072 0 1 1229
box 0 0 1 1
use contact_30  contact_30_527
timestamp 1634918361
transform 1 0 7072 0 1 1637
box 0 0 1 1
use contact_30  contact_30_528
timestamp 1634918361
transform 1 0 5304 0 1 31829
box 0 0 1 1
use contact_30  contact_30_529
timestamp 1634918361
transform 1 0 5304 0 1 31421
box 0 0 1 1
use contact_30  contact_30_530
timestamp 1634918361
transform 1 0 5440 0 1 1229
box 0 0 1 1
use contact_30  contact_30_531
timestamp 1634918361
transform 1 0 5440 0 1 1637
box 0 0 1 1
use contact_30  contact_30_532
timestamp 1634918361
transform 1 0 3808 0 1 1229
box 0 0 1 1
use contact_30  contact_30_533
timestamp 1634918361
transform 1 0 3808 0 1 1637
box 0 0 1 1
use contact_30  contact_30_534
timestamp 1634918361
transform 1 0 3808 0 1 31829
box 0 0 1 1
use contact_30  contact_30_535
timestamp 1634918361
transform 1 0 3808 0 1 31421
box 0 0 1 1
use contact_30  contact_30_536
timestamp 1634918361
transform 1 0 2176 0 1 31829
box 0 0 1 1
use contact_30  contact_30_537
timestamp 1634918361
transform 1 0 2176 0 1 31421
box 0 0 1 1
use contact_30  contact_30_538
timestamp 1634918361
transform 1 0 2176 0 1 1229
box 0 0 1 1
use contact_30  contact_30_539
timestamp 1634918361
transform 1 0 2176 0 1 1637
box 0 0 1 1
use contact_30  contact_30_540
timestamp 1634918361
transform 1 0 1224 0 1 23805
box 0 0 1 1
use contact_30  contact_30_541
timestamp 1634918361
transform 1 0 1224 0 1 10341
box 0 0 1 1
use contact_30  contact_30_542
timestamp 1634918361
transform 1 0 3264 0 1 11021
box 0 0 1 1
use contact_30  contact_30_543
timestamp 1634918361
transform 1 0 3264 0 1 10477
box 0 0 1 1
use contact_30  contact_30_544
timestamp 1634918361
transform 1 0 1224 0 1 15509
box 0 0 1 1
use contact_30  contact_30_545
timestamp 1634918361
transform 1 0 1224 0 1 8845
box 0 0 1 1
use contact_30  contact_30_546
timestamp 1634918361
transform 1 0 3264 0 1 8301
box 0 0 1 1
use contact_30  contact_30_547
timestamp 1634918361
transform 1 0 3264 0 1 8709
box 0 0 1 1
use contact_30  contact_30_548
timestamp 1634918361
transform 1 0 1224 0 1 27341
box 0 0 1 1
use contact_30  contact_30_549
timestamp 1634918361
transform 1 0 1224 0 1 13741
box 0 0 1 1
use contact_30  contact_30_550
timestamp 1634918361
transform 1 0 1224 0 1 7077
box 0 0 1 1
use contact_30  contact_30_551
timestamp 1634918361
transform 1 0 1224 0 1 17141
box 0 0 1 1
use contact_30  contact_30_552
timestamp 1634918361
transform 1 0 3264 0 1 16733
box 0 0 1 1
use contact_30  contact_30_553
timestamp 1634918361
transform 1 0 3264 0 1 17141
box 0 0 1 1
use contact_30  contact_30_554
timestamp 1634918361
transform 1 0 1224 0 1 25573
box 0 0 1 1
use contact_30  contact_30_555
timestamp 1634918361
transform 1 0 1224 0 1 12245
box 0 0 1 1
use contact_30  contact_30_556
timestamp 1634918361
transform 1 0 1224 0 1 20405
box 0 0 1 1
use contact_30  contact_30_557
timestamp 1634918361
transform 1 0 1224 0 1 28837
box 0 0 1 1
use contact_30  contact_30_558
timestamp 1634918361
transform 1 0 1224 0 1 30741
box 0 0 1 1
use contact_30  contact_30_559
timestamp 1634918361
transform 1 0 1224 0 1 18909
box 0 0 1 1
use contact_30  contact_30_560
timestamp 1634918361
transform 1 0 2448 0 1 19453
box 0 0 1 1
use contact_30  contact_30_561
timestamp 1634918361
transform 1 0 2448 0 1 18909
box 0 0 1 1
use contact_30  contact_30_562
timestamp 1634918361
transform 1 0 1224 0 1 5309
box 0 0 1 1
use contact_30  contact_30_563
timestamp 1634918361
transform 1 0 1224 0 1 22173
box 0 0 1 1
use contact_30  contact_30_564
timestamp 1634918361
transform 1 0 1224 0 1 3813
box 0 0 1 1
use contact_30  contact_30_565
timestamp 1634918361
transform 1 0 2040 0 1 1773
box 0 0 1 1
use contact_30  contact_30_566
timestamp 1634918361
transform 1 0 2040 0 1 2045
box 0 0 1 1
use contact_36  contact_36_0
timestamp 1634918361
transform 1 0 42840 0 1 413
box 0 0 1 1
use contact_36  contact_36_1
timestamp 1634918361
transform 1 0 544 0 1 32781
box 0 0 1 1
use contact_36  contact_36_2
timestamp 1634918361
transform 1 0 408 0 1 32781
box 0 0 1 1
use contact_36  contact_36_3
timestamp 1634918361
transform 1 0 272 0 1 549
box 0 0 1 1
use contact_36  contact_36_4
timestamp 1634918361
transform 1 0 42840 0 1 32509
box 0 0 1 1
use contact_36  contact_36_5
timestamp 1634918361
transform 1 0 272 0 1 277
box 0 0 1 1
use contact_36  contact_36_6
timestamp 1634918361
transform 1 0 43112 0 1 413
box 0 0 1 1
use contact_36  contact_36_7
timestamp 1634918361
transform 1 0 544 0 1 32509
box 0 0 1 1
use contact_36  contact_36_8
timestamp 1634918361
transform 1 0 42840 0 1 32781
box 0 0 1 1
use contact_36  contact_36_9
timestamp 1634918361
transform 1 0 42976 0 1 413
box 0 0 1 1
use contact_36  contact_36_10
timestamp 1634918361
transform 1 0 272 0 1 32645
box 0 0 1 1
use contact_36  contact_36_11
timestamp 1634918361
transform 1 0 408 0 1 32509
box 0 0 1 1
use contact_36  contact_36_12
timestamp 1634918361
transform 1 0 408 0 1 549
box 0 0 1 1
use contact_36  contact_36_13
timestamp 1634918361
transform 1 0 42840 0 1 277
box 0 0 1 1
use contact_36  contact_36_14
timestamp 1634918361
transform 1 0 43112 0 1 32781
box 0 0 1 1
use contact_36  contact_36_15
timestamp 1634918361
transform 1 0 544 0 1 549
box 0 0 1 1
use contact_36  contact_36_16
timestamp 1634918361
transform 1 0 42976 0 1 32781
box 0 0 1 1
use contact_36  contact_36_17
timestamp 1634918361
transform 1 0 544 0 1 277
box 0 0 1 1
use contact_36  contact_36_18
timestamp 1634918361
transform 1 0 42840 0 1 549
box 0 0 1 1
use contact_36  contact_36_19
timestamp 1634918361
transform 1 0 42976 0 1 32509
box 0 0 1 1
use contact_36  contact_36_20
timestamp 1634918361
transform 1 0 272 0 1 413
box 0 0 1 1
use contact_36  contact_36_21
timestamp 1634918361
transform 1 0 544 0 1 32645
box 0 0 1 1
use contact_36  contact_36_22
timestamp 1634918361
transform 1 0 43112 0 1 32509
box 0 0 1 1
use contact_36  contact_36_23
timestamp 1634918361
transform 1 0 408 0 1 277
box 0 0 1 1
use contact_36  contact_36_24
timestamp 1634918361
transform 1 0 42840 0 1 32645
box 0 0 1 1
use contact_36  contact_36_25
timestamp 1634918361
transform 1 0 408 0 1 32645
box 0 0 1 1
use contact_36  contact_36_26
timestamp 1634918361
transform 1 0 42976 0 1 549
box 0 0 1 1
use contact_36  contact_36_27
timestamp 1634918361
transform 1 0 272 0 1 32781
box 0 0 1 1
use contact_36  contact_36_28
timestamp 1634918361
transform 1 0 42976 0 1 277
box 0 0 1 1
use contact_36  contact_36_29
timestamp 1634918361
transform 1 0 43112 0 1 549
box 0 0 1 1
use contact_36  contact_36_30
timestamp 1634918361
transform 1 0 544 0 1 413
box 0 0 1 1
use contact_36  contact_36_31
timestamp 1634918361
transform 1 0 43112 0 1 277
box 0 0 1 1
use contact_36  contact_36_32
timestamp 1634918361
transform 1 0 408 0 1 413
box 0 0 1 1
use contact_36  contact_36_33
timestamp 1634918361
transform 1 0 272 0 1 32509
box 0 0 1 1
use contact_36  contact_36_34
timestamp 1634918361
transform 1 0 43112 0 1 32645
box 0 0 1 1
use contact_36  contact_36_35
timestamp 1634918361
transform 1 0 42976 0 1 32645
box 0 0 1 1
use contact_36  contact_36_36
timestamp 1634918361
transform 1 0 952 0 1 957
box 0 0 1 1
use contact_36  contact_36_37
timestamp 1634918361
transform 1 0 952 0 1 32101
box 0 0 1 1
use contact_36  contact_36_38
timestamp 1634918361
transform 1 0 42296 0 1 1093
box 0 0 1 1
use contact_36  contact_36_39
timestamp 1634918361
transform 1 0 42432 0 1 31965
box 0 0 1 1
use contact_36  contact_36_40
timestamp 1634918361
transform 1 0 42296 0 1 31965
box 0 0 1 1
use contact_36  contact_36_41
timestamp 1634918361
transform 1 0 42160 0 1 1229
box 0 0 1 1
use contact_36  contact_36_42
timestamp 1634918361
transform 1 0 1088 0 1 1229
box 0 0 1 1
use contact_36  contact_36_43
timestamp 1634918361
transform 1 0 42160 0 1 957
box 0 0 1 1
use contact_36  contact_36_44
timestamp 1634918361
transform 1 0 952 0 1 31829
box 0 0 1 1
use contact_36  contact_36_45
timestamp 1634918361
transform 1 0 1088 0 1 957
box 0 0 1 1
use contact_36  contact_36_46
timestamp 1634918361
transform 1 0 1224 0 1 1229
box 0 0 1 1
use contact_36  contact_36_47
timestamp 1634918361
transform 1 0 1224 0 1 957
box 0 0 1 1
use contact_36  contact_36_48
timestamp 1634918361
transform 1 0 952 0 1 1093
box 0 0 1 1
use contact_36  contact_36_49
timestamp 1634918361
transform 1 0 1224 0 1 32101
box 0 0 1 1
use contact_36  contact_36_50
timestamp 1634918361
transform 1 0 42160 0 1 32101
box 0 0 1 1
use contact_36  contact_36_51
timestamp 1634918361
transform 1 0 1224 0 1 31829
box 0 0 1 1
use contact_36  contact_36_52
timestamp 1634918361
transform 1 0 42296 0 1 1229
box 0 0 1 1
use contact_36  contact_36_53
timestamp 1634918361
transform 1 0 1088 0 1 32101
box 0 0 1 1
use contact_36  contact_36_54
timestamp 1634918361
transform 1 0 42160 0 1 31829
box 0 0 1 1
use contact_36  contact_36_55
timestamp 1634918361
transform 1 0 42296 0 1 957
box 0 0 1 1
use contact_36  contact_36_56
timestamp 1634918361
transform 1 0 42432 0 1 1093
box 0 0 1 1
use contact_36  contact_36_57
timestamp 1634918361
transform 1 0 1088 0 1 31829
box 0 0 1 1
use contact_36  contact_36_58
timestamp 1634918361
transform 1 0 42432 0 1 1229
box 0 0 1 1
use contact_36  contact_36_59
timestamp 1634918361
transform 1 0 42432 0 1 957
box 0 0 1 1
use contact_36  contact_36_60
timestamp 1634918361
transform 1 0 952 0 1 31965
box 0 0 1 1
use contact_36  contact_36_61
timestamp 1634918361
transform 1 0 42296 0 1 32101
box 0 0 1 1
use contact_36  contact_36_62
timestamp 1634918361
transform 1 0 1224 0 1 1093
box 0 0 1 1
use contact_36  contact_36_63
timestamp 1634918361
transform 1 0 42296 0 1 31829
box 0 0 1 1
use contact_36  contact_36_64
timestamp 1634918361
transform 1 0 42160 0 1 1093
box 0 0 1 1
use contact_36  contact_36_65
timestamp 1634918361
transform 1 0 42432 0 1 32101
box 0 0 1 1
use contact_36  contact_36_66
timestamp 1634918361
transform 1 0 1088 0 1 1093
box 0 0 1 1
use contact_36  contact_36_67
timestamp 1634918361
transform 1 0 42432 0 1 31829
box 0 0 1 1
use contact_36  contact_36_68
timestamp 1634918361
transform 1 0 42160 0 1 31965
box 0 0 1 1
use contact_36  contact_36_69
timestamp 1634918361
transform 1 0 1088 0 1 31965
box 0 0 1 1
use contact_36  contact_36_70
timestamp 1634918361
transform 1 0 1224 0 1 31965
box 0 0 1 1
use contact_36  contact_36_71
timestamp 1634918361
transform 1 0 952 0 1 1229
box 0 0 1 1
use contact_30  contact_30_567
timestamp 1634918361
transform 1 0 24072 0 1 10477
box 0 0 1 1
use contact_30  contact_30_568
timestamp 1634918361
transform 1 0 23664 0 1 10749
box 0 0 1 1
use contact_30  contact_30_569
timestamp 1634918361
transform 1 0 22848 0 1 10477
box 0 0 1 1
use contact_30  contact_30_570
timestamp 1634918361
transform 1 0 22440 0 1 10749
box 0 0 1 1
use contact_30  contact_30_571
timestamp 1634918361
transform 1 0 21624 0 1 10477
box 0 0 1 1
use contact_30  contact_30_572
timestamp 1634918361
transform 1 0 20944 0 1 10749
box 0 0 1 1
use contact_30  contact_30_573
timestamp 1634918361
transform 1 0 20264 0 1 10477
box 0 0 1 1
use contact_30  contact_30_574
timestamp 1634918361
transform 1 0 19720 0 1 10749
box 0 0 1 1
use contact_30  contact_30_575
timestamp 1634918361
transform 1 0 24208 0 1 25437
box 0 0 1 1
use contact_30  contact_30_576
timestamp 1634918361
transform 1 0 23120 0 1 25437
box 0 0 1 1
use contact_30  contact_30_577
timestamp 1634918361
transform 1 0 22848 0 1 25437
box 0 0 1 1
use contact_30  contact_30_578
timestamp 1634918361
transform 1 0 21896 0 1 25437
box 0 0 1 1
use contact_30  contact_30_579
timestamp 1634918361
transform 1 0 21624 0 1 25437
box 0 0 1 1
use contact_30  contact_30_580
timestamp 1634918361
transform 1 0 20672 0 1 25437
box 0 0 1 1
use contact_30  contact_30_581
timestamp 1634918361
transform 1 0 20400 0 1 25437
box 0 0 1 1
use contact_30  contact_30_582
timestamp 1634918361
transform 1 0 19312 0 1 25437
box 0 0 1 1
use contact_30  contact_30_583
timestamp 1634918361
transform 1 0 8568 0 1 26253
box 0 0 1 1
use contact_30  contact_30_584
timestamp 1634918361
transform 1 0 37400 0 1 29925
box 0 0 1 1
use contact_30  contact_30_585
timestamp 1634918361
transform 1 0 5984 0 1 3133
box 0 0 1 1
use contact_30  contact_30_586
timestamp 1634918361
transform 1 0 14416 0 1 3133
box 0 0 1 1
use contact_30  contact_30_587
timestamp 1634918361
transform 1 0 13192 0 1 3133
box 0 0 1 1
use contact_30  contact_30_588
timestamp 1634918361
transform 1 0 12104 0 1 3133
box 0 0 1 1
use contact_30  contact_30_589
timestamp 1634918361
transform 1 0 10744 0 1 3133
box 0 0 1 1
use contact_30  contact_30_590
timestamp 1634918361
transform 1 0 23800 0 1 3133
box 0 0 1 1
use contact_30  contact_30_591
timestamp 1634918361
transform 1 0 22576 0 1 3133
box 0 0 1 1
use contact_30  contact_30_592
timestamp 1634918361
transform 1 0 21352 0 1 3133
box 0 0 1 1
use contact_30  contact_30_593
timestamp 1634918361
transform 1 0 20264 0 1 3133
box 0 0 1 1
use contact_30  contact_30_594
timestamp 1634918361
transform 1 0 19040 0 1 3133
box 0 0 1 1
use contact_30  contact_30_595
timestamp 1634918361
transform 1 0 17952 0 1 3133
box 0 0 1 1
use contact_30  contact_30_596
timestamp 1634918361
transform 1 0 16728 0 1 3133
box 0 0 1 1
use contact_30  contact_30_597
timestamp 1634918361
transform 1 0 15504 0 1 3133
box 0 0 1 1
use contact_35  contact_35_0
timestamp 1634918361
transform 1 0 1662 0 1 31288
box 0 0 192 192
use contact_35  contact_35_1
timestamp 1634918361
transform 1 0 41644 0 1 31288
box 0 0 192 192
use contact_35  contact_35_2
timestamp 1634918361
transform 1 0 41644 0 1 1664
box 0 0 192 192
use contact_35  contact_35_3
timestamp 1634918361
transform 1 0 1662 0 1 1664
box 0 0 192 192
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 41708 0 1 30960
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1634918361
transform 1 0 41711 0 1 30959
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1634918361
transform 1 0 41715 0 1 30951
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 41707 0 1 30619
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 41708 0 1 30624
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1634918361
transform 1 0 41711 0 1 30623
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1634918361
transform 1 0 41715 0 1 30615
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 41708 0 1 30288
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1634918361
transform 1 0 41711 0 1 30287
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1634918361
transform 1 0 41715 0 1 30279
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 41708 0 1 29952
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1634918361
transform 1 0 41711 0 1 29951
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1634918361
transform 1 0 41715 0 1 29943
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 41708 0 1 29616
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1634918361
transform 1 0 41711 0 1 29615
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1634918361
transform 1 0 41715 0 1 29607
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 41708 0 1 29280
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1634918361
transform 1 0 41711 0 1 29279
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1634918361
transform 1 0 41715 0 1 29271
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 41707 0 1 28939
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 41708 0 1 28944
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1634918361
transform 1 0 41711 0 1 28943
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1634918361
transform 1 0 41715 0 1 28935
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 41708 0 1 28608
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1634918361
transform 1 0 41711 0 1 28607
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1634918361
transform 1 0 41715 0 1 28599
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1634918361
transform 1 0 41708 0 1 28272
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1634918361
transform 1 0 41711 0 1 28271
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1634918361
transform 1 0 41715 0 1 28263
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1634918361
transform 1 0 41708 0 1 27936
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1634918361
transform 1 0 41711 0 1 27935
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1634918361
transform 1 0 41715 0 1 27927
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1634918361
transform 1 0 41708 0 1 27600
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1634918361
transform 1 0 41711 0 1 27599
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1634918361
transform 1 0 41715 0 1 27591
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 41707 0 1 27259
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1634918361
transform 1 0 41708 0 1 27264
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1634918361
transform 1 0 41711 0 1 27263
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1634918361
transform 1 0 41715 0 1 27255
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1634918361
transform 1 0 41708 0 1 26928
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1634918361
transform 1 0 41711 0 1 26927
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1634918361
transform 1 0 41715 0 1 26919
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1634918361
transform 1 0 41708 0 1 26592
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1634918361
transform 1 0 41711 0 1 26591
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1634918361
transform 1 0 41715 0 1 26583
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1634918361
transform 1 0 41708 0 1 26256
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1634918361
transform 1 0 41711 0 1 26255
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1634918361
transform 1 0 41715 0 1 26247
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1634918361
transform 1 0 41708 0 1 25920
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1634918361
transform 1 0 41711 0 1 25919
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1634918361
transform 1 0 41715 0 1 25911
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 41707 0 1 25579
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1634918361
transform 1 0 41708 0 1 25584
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1634918361
transform 1 0 41711 0 1 25583
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1634918361
transform 1 0 41715 0 1 25575
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1634918361
transform 1 0 41708 0 1 25248
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1634918361
transform 1 0 41711 0 1 25247
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1634918361
transform 1 0 41715 0 1 25239
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1634918361
transform 1 0 41708 0 1 24912
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1634918361
transform 1 0 41711 0 1 24911
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1634918361
transform 1 0 41715 0 1 24903
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1634918361
transform 1 0 41708 0 1 24576
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1634918361
transform 1 0 41711 0 1 24575
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1634918361
transform 1 0 41715 0 1 24567
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1634918361
transform 1 0 41708 0 1 24240
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1634918361
transform 1 0 41711 0 1 24239
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1634918361
transform 1 0 41715 0 1 24231
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 41707 0 1 23899
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1634918361
transform 1 0 41708 0 1 23904
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1634918361
transform 1 0 41711 0 1 23903
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1634918361
transform 1 0 41715 0 1 23895
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1634918361
transform 1 0 41708 0 1 23568
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1634918361
transform 1 0 41711 0 1 23567
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1634918361
transform 1 0 41715 0 1 23559
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1634918361
transform 1 0 41708 0 1 23232
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1634918361
transform 1 0 41711 0 1 23231
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1634918361
transform 1 0 41715 0 1 23223
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1634918361
transform 1 0 41708 0 1 22896
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1634918361
transform 1 0 41711 0 1 22895
box 0 0 1 1
use contact_13  contact_13_24
timestamp 1634918361
transform 1 0 41715 0 1 22887
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1634918361
transform 1 0 41708 0 1 22560
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1634918361
transform 1 0 41711 0 1 22559
box 0 0 1 1
use contact_13  contact_13_25
timestamp 1634918361
transform 1 0 41715 0 1 22551
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 41707 0 1 22219
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1634918361
transform 1 0 41708 0 1 22224
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1634918361
transform 1 0 41711 0 1 22223
box 0 0 1 1
use contact_13  contact_13_26
timestamp 1634918361
transform 1 0 41715 0 1 22215
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1634918361
transform 1 0 41708 0 1 21888
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1634918361
transform 1 0 41711 0 1 21887
box 0 0 1 1
use contact_13  contact_13_27
timestamp 1634918361
transform 1 0 41715 0 1 21879
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1634918361
transform 1 0 41708 0 1 21552
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1634918361
transform 1 0 41711 0 1 21551
box 0 0 1 1
use contact_13  contact_13_28
timestamp 1634918361
transform 1 0 41715 0 1 21543
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1634918361
transform 1 0 41708 0 1 21216
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1634918361
transform 1 0 41711 0 1 21215
box 0 0 1 1
use contact_13  contact_13_29
timestamp 1634918361
transform 1 0 41715 0 1 21207
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1634918361
transform 1 0 41708 0 1 20880
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1634918361
transform 1 0 41711 0 1 20879
box 0 0 1 1
use contact_13  contact_13_30
timestamp 1634918361
transform 1 0 41715 0 1 20871
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 41707 0 1 20539
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1634918361
transform 1 0 41708 0 1 20544
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1634918361
transform 1 0 41711 0 1 20543
box 0 0 1 1
use contact_13  contact_13_31
timestamp 1634918361
transform 1 0 41715 0 1 20535
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1634918361
transform 1 0 41708 0 1 20208
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1634918361
transform 1 0 41711 0 1 20207
box 0 0 1 1
use contact_13  contact_13_32
timestamp 1634918361
transform 1 0 41715 0 1 20199
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1634918361
transform 1 0 41708 0 1 19872
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1634918361
transform 1 0 41711 0 1 19871
box 0 0 1 1
use contact_13  contact_13_33
timestamp 1634918361
transform 1 0 41715 0 1 19863
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1634918361
transform 1 0 41708 0 1 19536
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1634918361
transform 1 0 41711 0 1 19535
box 0 0 1 1
use contact_13  contact_13_34
timestamp 1634918361
transform 1 0 41715 0 1 19527
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1634918361
transform 1 0 41708 0 1 19200
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1634918361
transform 1 0 41711 0 1 19199
box 0 0 1 1
use contact_13  contact_13_35
timestamp 1634918361
transform 1 0 41715 0 1 19191
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 41707 0 1 18859
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1634918361
transform 1 0 41708 0 1 18864
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1634918361
transform 1 0 41711 0 1 18863
box 0 0 1 1
use contact_13  contact_13_36
timestamp 1634918361
transform 1 0 41715 0 1 18855
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1634918361
transform 1 0 41708 0 1 18528
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1634918361
transform 1 0 41711 0 1 18527
box 0 0 1 1
use contact_13  contact_13_37
timestamp 1634918361
transform 1 0 41715 0 1 18519
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1634918361
transform 1 0 41708 0 1 18192
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1634918361
transform 1 0 41711 0 1 18191
box 0 0 1 1
use contact_13  contact_13_38
timestamp 1634918361
transform 1 0 41715 0 1 18183
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1634918361
transform 1 0 41708 0 1 17856
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1634918361
transform 1 0 41711 0 1 17855
box 0 0 1 1
use contact_13  contact_13_39
timestamp 1634918361
transform 1 0 41715 0 1 17847
box 0 0 1 1
use contact_19  contact_19_40
timestamp 1634918361
transform 1 0 41708 0 1 17520
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1634918361
transform 1 0 41711 0 1 17519
box 0 0 1 1
use contact_13  contact_13_40
timestamp 1634918361
transform 1 0 41715 0 1 17511
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 41707 0 1 17179
box 0 0 1 1
use contact_19  contact_19_41
timestamp 1634918361
transform 1 0 41708 0 1 17184
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1634918361
transform 1 0 41711 0 1 17183
box 0 0 1 1
use contact_13  contact_13_41
timestamp 1634918361
transform 1 0 41715 0 1 17175
box 0 0 1 1
use contact_19  contact_19_42
timestamp 1634918361
transform 1 0 41708 0 1 16848
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1634918361
transform 1 0 41711 0 1 16847
box 0 0 1 1
use contact_13  contact_13_42
timestamp 1634918361
transform 1 0 41715 0 1 16839
box 0 0 1 1
use contact_19  contact_19_43
timestamp 1634918361
transform 1 0 41708 0 1 16512
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1634918361
transform 1 0 41711 0 1 16511
box 0 0 1 1
use contact_13  contact_13_43
timestamp 1634918361
transform 1 0 41715 0 1 16503
box 0 0 1 1
use contact_19  contact_19_44
timestamp 1634918361
transform 1 0 41708 0 1 16176
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1634918361
transform 1 0 41711 0 1 16175
box 0 0 1 1
use contact_13  contact_13_44
timestamp 1634918361
transform 1 0 41715 0 1 16167
box 0 0 1 1
use contact_19  contact_19_45
timestamp 1634918361
transform 1 0 41708 0 1 15840
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1634918361
transform 1 0 41711 0 1 15839
box 0 0 1 1
use contact_13  contact_13_45
timestamp 1634918361
transform 1 0 41715 0 1 15831
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 41707 0 1 15499
box 0 0 1 1
use contact_19  contact_19_46
timestamp 1634918361
transform 1 0 41708 0 1 15504
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1634918361
transform 1 0 41711 0 1 15503
box 0 0 1 1
use contact_13  contact_13_46
timestamp 1634918361
transform 1 0 41715 0 1 15495
box 0 0 1 1
use contact_19  contact_19_47
timestamp 1634918361
transform 1 0 41708 0 1 15168
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1634918361
transform 1 0 41711 0 1 15167
box 0 0 1 1
use contact_13  contact_13_47
timestamp 1634918361
transform 1 0 41715 0 1 15159
box 0 0 1 1
use contact_19  contact_19_48
timestamp 1634918361
transform 1 0 41708 0 1 14832
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1634918361
transform 1 0 41711 0 1 14831
box 0 0 1 1
use contact_13  contact_13_48
timestamp 1634918361
transform 1 0 41715 0 1 14823
box 0 0 1 1
use contact_19  contact_19_49
timestamp 1634918361
transform 1 0 41708 0 1 14496
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1634918361
transform 1 0 41711 0 1 14495
box 0 0 1 1
use contact_13  contact_13_49
timestamp 1634918361
transform 1 0 41715 0 1 14487
box 0 0 1 1
use contact_19  contact_19_50
timestamp 1634918361
transform 1 0 41708 0 1 14160
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1634918361
transform 1 0 41711 0 1 14159
box 0 0 1 1
use contact_13  contact_13_50
timestamp 1634918361
transform 1 0 41715 0 1 14151
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 41707 0 1 13819
box 0 0 1 1
use contact_19  contact_19_51
timestamp 1634918361
transform 1 0 41708 0 1 13824
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1634918361
transform 1 0 41711 0 1 13823
box 0 0 1 1
use contact_13  contact_13_51
timestamp 1634918361
transform 1 0 41715 0 1 13815
box 0 0 1 1
use contact_19  contact_19_52
timestamp 1634918361
transform 1 0 41708 0 1 13488
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1634918361
transform 1 0 41711 0 1 13487
box 0 0 1 1
use contact_13  contact_13_52
timestamp 1634918361
transform 1 0 41715 0 1 13479
box 0 0 1 1
use contact_19  contact_19_53
timestamp 1634918361
transform 1 0 41708 0 1 13152
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1634918361
transform 1 0 41711 0 1 13151
box 0 0 1 1
use contact_13  contact_13_53
timestamp 1634918361
transform 1 0 41715 0 1 13143
box 0 0 1 1
use contact_19  contact_19_54
timestamp 1634918361
transform 1 0 41708 0 1 12816
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1634918361
transform 1 0 41711 0 1 12815
box 0 0 1 1
use contact_13  contact_13_54
timestamp 1634918361
transform 1 0 41715 0 1 12807
box 0 0 1 1
use contact_19  contact_19_55
timestamp 1634918361
transform 1 0 41708 0 1 12480
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1634918361
transform 1 0 41711 0 1 12479
box 0 0 1 1
use contact_13  contact_13_55
timestamp 1634918361
transform 1 0 41715 0 1 12471
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 41707 0 1 12139
box 0 0 1 1
use contact_19  contact_19_56
timestamp 1634918361
transform 1 0 41708 0 1 12144
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1634918361
transform 1 0 41711 0 1 12143
box 0 0 1 1
use contact_13  contact_13_56
timestamp 1634918361
transform 1 0 41715 0 1 12135
box 0 0 1 1
use contact_19  contact_19_57
timestamp 1634918361
transform 1 0 41708 0 1 11808
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1634918361
transform 1 0 41711 0 1 11807
box 0 0 1 1
use contact_13  contact_13_57
timestamp 1634918361
transform 1 0 41715 0 1 11799
box 0 0 1 1
use contact_19  contact_19_58
timestamp 1634918361
transform 1 0 41708 0 1 11472
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1634918361
transform 1 0 41711 0 1 11471
box 0 0 1 1
use contact_13  contact_13_58
timestamp 1634918361
transform 1 0 41715 0 1 11463
box 0 0 1 1
use contact_19  contact_19_59
timestamp 1634918361
transform 1 0 41708 0 1 11136
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1634918361
transform 1 0 41711 0 1 11135
box 0 0 1 1
use contact_13  contact_13_59
timestamp 1634918361
transform 1 0 41715 0 1 11127
box 0 0 1 1
use contact_19  contact_19_60
timestamp 1634918361
transform 1 0 41708 0 1 10800
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1634918361
transform 1 0 41711 0 1 10799
box 0 0 1 1
use contact_13  contact_13_60
timestamp 1634918361
transform 1 0 41715 0 1 10791
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 41707 0 1 10459
box 0 0 1 1
use contact_19  contact_19_61
timestamp 1634918361
transform 1 0 41708 0 1 10464
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1634918361
transform 1 0 41711 0 1 10463
box 0 0 1 1
use contact_13  contact_13_61
timestamp 1634918361
transform 1 0 41715 0 1 10455
box 0 0 1 1
use contact_19  contact_19_62
timestamp 1634918361
transform 1 0 41708 0 1 10128
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1634918361
transform 1 0 41711 0 1 10127
box 0 0 1 1
use contact_13  contact_13_62
timestamp 1634918361
transform 1 0 41715 0 1 10119
box 0 0 1 1
use contact_19  contact_19_63
timestamp 1634918361
transform 1 0 41708 0 1 9792
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1634918361
transform 1 0 41711 0 1 9791
box 0 0 1 1
use contact_13  contact_13_63
timestamp 1634918361
transform 1 0 41715 0 1 9783
box 0 0 1 1
use contact_19  contact_19_64
timestamp 1634918361
transform 1 0 41708 0 1 9456
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1634918361
transform 1 0 41711 0 1 9455
box 0 0 1 1
use contact_13  contact_13_64
timestamp 1634918361
transform 1 0 41715 0 1 9447
box 0 0 1 1
use contact_19  contact_19_65
timestamp 1634918361
transform 1 0 41708 0 1 9120
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1634918361
transform 1 0 41711 0 1 9119
box 0 0 1 1
use contact_13  contact_13_65
timestamp 1634918361
transform 1 0 41715 0 1 9111
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 41707 0 1 8779
box 0 0 1 1
use contact_19  contact_19_66
timestamp 1634918361
transform 1 0 41708 0 1 8784
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1634918361
transform 1 0 41711 0 1 8783
box 0 0 1 1
use contact_13  contact_13_66
timestamp 1634918361
transform 1 0 41715 0 1 8775
box 0 0 1 1
use contact_19  contact_19_67
timestamp 1634918361
transform 1 0 41708 0 1 8448
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1634918361
transform 1 0 41711 0 1 8447
box 0 0 1 1
use contact_13  contact_13_67
timestamp 1634918361
transform 1 0 41715 0 1 8439
box 0 0 1 1
use contact_19  contact_19_68
timestamp 1634918361
transform 1 0 41708 0 1 8112
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1634918361
transform 1 0 41711 0 1 8111
box 0 0 1 1
use contact_13  contact_13_68
timestamp 1634918361
transform 1 0 41715 0 1 8103
box 0 0 1 1
use contact_19  contact_19_69
timestamp 1634918361
transform 1 0 41708 0 1 7776
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1634918361
transform 1 0 41711 0 1 7775
box 0 0 1 1
use contact_13  contact_13_69
timestamp 1634918361
transform 1 0 41715 0 1 7767
box 0 0 1 1
use contact_19  contact_19_70
timestamp 1634918361
transform 1 0 41708 0 1 7440
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1634918361
transform 1 0 41711 0 1 7439
box 0 0 1 1
use contact_13  contact_13_70
timestamp 1634918361
transform 1 0 41715 0 1 7431
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 41707 0 1 7099
box 0 0 1 1
use contact_19  contact_19_71
timestamp 1634918361
transform 1 0 41708 0 1 7104
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1634918361
transform 1 0 41711 0 1 7103
box 0 0 1 1
use contact_13  contact_13_71
timestamp 1634918361
transform 1 0 41715 0 1 7095
box 0 0 1 1
use contact_19  contact_19_72
timestamp 1634918361
transform 1 0 41708 0 1 6768
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1634918361
transform 1 0 41711 0 1 6767
box 0 0 1 1
use contact_13  contact_13_72
timestamp 1634918361
transform 1 0 41715 0 1 6759
box 0 0 1 1
use contact_19  contact_19_73
timestamp 1634918361
transform 1 0 41708 0 1 6432
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1634918361
transform 1 0 41711 0 1 6431
box 0 0 1 1
use contact_13  contact_13_73
timestamp 1634918361
transform 1 0 41715 0 1 6423
box 0 0 1 1
use contact_19  contact_19_74
timestamp 1634918361
transform 1 0 41708 0 1 6096
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1634918361
transform 1 0 41711 0 1 6095
box 0 0 1 1
use contact_13  contact_13_74
timestamp 1634918361
transform 1 0 41715 0 1 6087
box 0 0 1 1
use contact_19  contact_19_75
timestamp 1634918361
transform 1 0 41708 0 1 5760
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1634918361
transform 1 0 41711 0 1 5759
box 0 0 1 1
use contact_13  contact_13_75
timestamp 1634918361
transform 1 0 41715 0 1 5751
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 41707 0 1 5419
box 0 0 1 1
use contact_19  contact_19_76
timestamp 1634918361
transform 1 0 41708 0 1 5424
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1634918361
transform 1 0 41711 0 1 5423
box 0 0 1 1
use contact_13  contact_13_76
timestamp 1634918361
transform 1 0 41715 0 1 5415
box 0 0 1 1
use contact_19  contact_19_77
timestamp 1634918361
transform 1 0 41708 0 1 5088
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1634918361
transform 1 0 41711 0 1 5087
box 0 0 1 1
use contact_13  contact_13_77
timestamp 1634918361
transform 1 0 41715 0 1 5079
box 0 0 1 1
use contact_19  contact_19_78
timestamp 1634918361
transform 1 0 41708 0 1 4752
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1634918361
transform 1 0 41711 0 1 4751
box 0 0 1 1
use contact_13  contact_13_78
timestamp 1634918361
transform 1 0 41715 0 1 4743
box 0 0 1 1
use contact_19  contact_19_79
timestamp 1634918361
transform 1 0 41708 0 1 4416
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1634918361
transform 1 0 41711 0 1 4415
box 0 0 1 1
use contact_13  contact_13_79
timestamp 1634918361
transform 1 0 41715 0 1 4407
box 0 0 1 1
use contact_19  contact_19_80
timestamp 1634918361
transform 1 0 41708 0 1 4080
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1634918361
transform 1 0 41711 0 1 4079
box 0 0 1 1
use contact_13  contact_13_80
timestamp 1634918361
transform 1 0 41715 0 1 4071
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 41707 0 1 3739
box 0 0 1 1
use contact_19  contact_19_81
timestamp 1634918361
transform 1 0 41708 0 1 3744
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1634918361
transform 1 0 41711 0 1 3743
box 0 0 1 1
use contact_13  contact_13_81
timestamp 1634918361
transform 1 0 41715 0 1 3735
box 0 0 1 1
use contact_19  contact_19_82
timestamp 1634918361
transform 1 0 41708 0 1 3408
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1634918361
transform 1 0 41711 0 1 3407
box 0 0 1 1
use contact_13  contact_13_82
timestamp 1634918361
transform 1 0 41715 0 1 3399
box 0 0 1 1
use contact_19  contact_19_83
timestamp 1634918361
transform 1 0 41708 0 1 3072
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1634918361
transform 1 0 41711 0 1 3071
box 0 0 1 1
use contact_13  contact_13_83
timestamp 1634918361
transform 1 0 41715 0 1 3063
box 0 0 1 1
use contact_19  contact_19_84
timestamp 1634918361
transform 1 0 41708 0 1 2736
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1634918361
transform 1 0 41711 0 1 2735
box 0 0 1 1
use contact_13  contact_13_84
timestamp 1634918361
transform 1 0 41715 0 1 2727
box 0 0 1 1
use contact_19  contact_19_85
timestamp 1634918361
transform 1 0 41708 0 1 2400
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1634918361
transform 1 0 41711 0 1 2399
box 0 0 1 1
use contact_13  contact_13_85
timestamp 1634918361
transform 1 0 41715 0 1 2391
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1634918361
transform 1 0 41707 0 1 2059
box 0 0 1 1
use contact_19  contact_19_86
timestamp 1634918361
transform 1 0 41708 0 1 2064
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1634918361
transform 1 0 41711 0 1 2063
box 0 0 1 1
use contact_13  contact_13_86
timestamp 1634918361
transform 1 0 41715 0 1 2055
box 0 0 1 1
use contact_19  contact_19_87
timestamp 1634918361
transform 1 0 1726 0 1 30960
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1634918361
transform 1 0 1729 0 1 30959
box 0 0 1 1
use contact_13  contact_13_87
timestamp 1634918361
transform 1 0 1733 0 1 30951
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1634918361
transform 1 0 1725 0 1 30619
box 0 0 1 1
use contact_19  contact_19_88
timestamp 1634918361
transform 1 0 1726 0 1 30624
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1634918361
transform 1 0 1729 0 1 30623
box 0 0 1 1
use contact_13  contact_13_88
timestamp 1634918361
transform 1 0 1733 0 1 30615
box 0 0 1 1
use contact_19  contact_19_89
timestamp 1634918361
transform 1 0 1726 0 1 30288
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1634918361
transform 1 0 1729 0 1 30287
box 0 0 1 1
use contact_13  contact_13_89
timestamp 1634918361
transform 1 0 1733 0 1 30279
box 0 0 1 1
use contact_19  contact_19_90
timestamp 1634918361
transform 1 0 1726 0 1 29952
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1634918361
transform 1 0 1729 0 1 29951
box 0 0 1 1
use contact_13  contact_13_90
timestamp 1634918361
transform 1 0 1733 0 1 29943
box 0 0 1 1
use contact_19  contact_19_91
timestamp 1634918361
transform 1 0 1726 0 1 29616
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1634918361
transform 1 0 1729 0 1 29615
box 0 0 1 1
use contact_13  contact_13_91
timestamp 1634918361
transform 1 0 1733 0 1 29607
box 0 0 1 1
use contact_19  contact_19_92
timestamp 1634918361
transform 1 0 1726 0 1 29280
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1634918361
transform 1 0 1729 0 1 29279
box 0 0 1 1
use contact_13  contact_13_92
timestamp 1634918361
transform 1 0 1733 0 1 29271
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1634918361
transform 1 0 1725 0 1 28939
box 0 0 1 1
use contact_19  contact_19_93
timestamp 1634918361
transform 1 0 1726 0 1 28944
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1634918361
transform 1 0 1729 0 1 28943
box 0 0 1 1
use contact_13  contact_13_93
timestamp 1634918361
transform 1 0 1733 0 1 28935
box 0 0 1 1
use contact_19  contact_19_94
timestamp 1634918361
transform 1 0 1726 0 1 28608
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1634918361
transform 1 0 1729 0 1 28607
box 0 0 1 1
use contact_13  contact_13_94
timestamp 1634918361
transform 1 0 1733 0 1 28599
box 0 0 1 1
use contact_19  contact_19_95
timestamp 1634918361
transform 1 0 1726 0 1 28272
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1634918361
transform 1 0 1729 0 1 28271
box 0 0 1 1
use contact_13  contact_13_95
timestamp 1634918361
transform 1 0 1733 0 1 28263
box 0 0 1 1
use contact_19  contact_19_96
timestamp 1634918361
transform 1 0 1726 0 1 27936
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1634918361
transform 1 0 1729 0 1 27935
box 0 0 1 1
use contact_13  contact_13_96
timestamp 1634918361
transform 1 0 1733 0 1 27927
box 0 0 1 1
use contact_19  contact_19_97
timestamp 1634918361
transform 1 0 1726 0 1 27600
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1634918361
transform 1 0 1729 0 1 27599
box 0 0 1 1
use contact_13  contact_13_97
timestamp 1634918361
transform 1 0 1733 0 1 27591
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1634918361
transform 1 0 1725 0 1 27259
box 0 0 1 1
use contact_19  contact_19_98
timestamp 1634918361
transform 1 0 1726 0 1 27264
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1634918361
transform 1 0 1729 0 1 27263
box 0 0 1 1
use contact_13  contact_13_98
timestamp 1634918361
transform 1 0 1733 0 1 27255
box 0 0 1 1
use contact_19  contact_19_99
timestamp 1634918361
transform 1 0 1726 0 1 26928
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1634918361
transform 1 0 1729 0 1 26927
box 0 0 1 1
use contact_13  contact_13_99
timestamp 1634918361
transform 1 0 1733 0 1 26919
box 0 0 1 1
use contact_19  contact_19_100
timestamp 1634918361
transform 1 0 1726 0 1 26592
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1634918361
transform 1 0 1729 0 1 26591
box 0 0 1 1
use contact_13  contact_13_100
timestamp 1634918361
transform 1 0 1733 0 1 26583
box 0 0 1 1
use contact_19  contact_19_101
timestamp 1634918361
transform 1 0 1726 0 1 26256
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1634918361
transform 1 0 1729 0 1 26255
box 0 0 1 1
use contact_13  contact_13_101
timestamp 1634918361
transform 1 0 1733 0 1 26247
box 0 0 1 1
use contact_19  contact_19_102
timestamp 1634918361
transform 1 0 1726 0 1 25920
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1634918361
transform 1 0 1729 0 1 25919
box 0 0 1 1
use contact_13  contact_13_102
timestamp 1634918361
transform 1 0 1733 0 1 25911
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1634918361
transform 1 0 1725 0 1 25579
box 0 0 1 1
use contact_19  contact_19_103
timestamp 1634918361
transform 1 0 1726 0 1 25584
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1634918361
transform 1 0 1729 0 1 25583
box 0 0 1 1
use contact_13  contact_13_103
timestamp 1634918361
transform 1 0 1733 0 1 25575
box 0 0 1 1
use contact_19  contact_19_104
timestamp 1634918361
transform 1 0 1726 0 1 25248
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1634918361
transform 1 0 1729 0 1 25247
box 0 0 1 1
use contact_13  contact_13_104
timestamp 1634918361
transform 1 0 1733 0 1 25239
box 0 0 1 1
use contact_19  contact_19_105
timestamp 1634918361
transform 1 0 1726 0 1 24912
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1634918361
transform 1 0 1729 0 1 24911
box 0 0 1 1
use contact_13  contact_13_105
timestamp 1634918361
transform 1 0 1733 0 1 24903
box 0 0 1 1
use contact_19  contact_19_106
timestamp 1634918361
transform 1 0 1726 0 1 24576
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1634918361
transform 1 0 1729 0 1 24575
box 0 0 1 1
use contact_13  contact_13_106
timestamp 1634918361
transform 1 0 1733 0 1 24567
box 0 0 1 1
use contact_19  contact_19_107
timestamp 1634918361
transform 1 0 1726 0 1 24240
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1634918361
transform 1 0 1729 0 1 24239
box 0 0 1 1
use contact_13  contact_13_107
timestamp 1634918361
transform 1 0 1733 0 1 24231
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1634918361
transform 1 0 1725 0 1 23899
box 0 0 1 1
use contact_19  contact_19_108
timestamp 1634918361
transform 1 0 1726 0 1 23904
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1634918361
transform 1 0 1729 0 1 23903
box 0 0 1 1
use contact_13  contact_13_108
timestamp 1634918361
transform 1 0 1733 0 1 23895
box 0 0 1 1
use contact_19  contact_19_109
timestamp 1634918361
transform 1 0 1726 0 1 23568
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1634918361
transform 1 0 1729 0 1 23567
box 0 0 1 1
use contact_13  contact_13_109
timestamp 1634918361
transform 1 0 1733 0 1 23559
box 0 0 1 1
use contact_19  contact_19_110
timestamp 1634918361
transform 1 0 1726 0 1 23232
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1634918361
transform 1 0 1729 0 1 23231
box 0 0 1 1
use contact_13  contact_13_110
timestamp 1634918361
transform 1 0 1733 0 1 23223
box 0 0 1 1
use contact_19  contact_19_111
timestamp 1634918361
transform 1 0 1726 0 1 22896
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1634918361
transform 1 0 1729 0 1 22895
box 0 0 1 1
use contact_13  contact_13_111
timestamp 1634918361
transform 1 0 1733 0 1 22887
box 0 0 1 1
use contact_19  contact_19_112
timestamp 1634918361
transform 1 0 1726 0 1 22560
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1634918361
transform 1 0 1729 0 1 22559
box 0 0 1 1
use contact_13  contact_13_112
timestamp 1634918361
transform 1 0 1733 0 1 22551
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1634918361
transform 1 0 1725 0 1 22219
box 0 0 1 1
use contact_19  contact_19_113
timestamp 1634918361
transform 1 0 1726 0 1 22224
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1634918361
transform 1 0 1729 0 1 22223
box 0 0 1 1
use contact_13  contact_13_113
timestamp 1634918361
transform 1 0 1733 0 1 22215
box 0 0 1 1
use contact_19  contact_19_114
timestamp 1634918361
transform 1 0 1726 0 1 21888
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1634918361
transform 1 0 1729 0 1 21887
box 0 0 1 1
use contact_13  contact_13_114
timestamp 1634918361
transform 1 0 1733 0 1 21879
box 0 0 1 1
use contact_19  contact_19_115
timestamp 1634918361
transform 1 0 1726 0 1 21552
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1634918361
transform 1 0 1729 0 1 21551
box 0 0 1 1
use contact_13  contact_13_115
timestamp 1634918361
transform 1 0 1733 0 1 21543
box 0 0 1 1
use contact_19  contact_19_116
timestamp 1634918361
transform 1 0 1726 0 1 21216
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1634918361
transform 1 0 1729 0 1 21215
box 0 0 1 1
use contact_13  contact_13_116
timestamp 1634918361
transform 1 0 1733 0 1 21207
box 0 0 1 1
use contact_19  contact_19_117
timestamp 1634918361
transform 1 0 1726 0 1 20880
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1634918361
transform 1 0 1729 0 1 20879
box 0 0 1 1
use contact_13  contact_13_117
timestamp 1634918361
transform 1 0 1733 0 1 20871
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1634918361
transform 1 0 1725 0 1 20539
box 0 0 1 1
use contact_19  contact_19_118
timestamp 1634918361
transform 1 0 1726 0 1 20544
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1634918361
transform 1 0 1729 0 1 20543
box 0 0 1 1
use contact_13  contact_13_118
timestamp 1634918361
transform 1 0 1733 0 1 20535
box 0 0 1 1
use contact_19  contact_19_119
timestamp 1634918361
transform 1 0 1726 0 1 20208
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1634918361
transform 1 0 1729 0 1 20207
box 0 0 1 1
use contact_13  contact_13_119
timestamp 1634918361
transform 1 0 1733 0 1 20199
box 0 0 1 1
use contact_19  contact_19_120
timestamp 1634918361
transform 1 0 1726 0 1 19872
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1634918361
transform 1 0 1729 0 1 19871
box 0 0 1 1
use contact_13  contact_13_120
timestamp 1634918361
transform 1 0 1733 0 1 19863
box 0 0 1 1
use contact_19  contact_19_121
timestamp 1634918361
transform 1 0 1726 0 1 19536
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1634918361
transform 1 0 1729 0 1 19535
box 0 0 1 1
use contact_13  contact_13_121
timestamp 1634918361
transform 1 0 1733 0 1 19527
box 0 0 1 1
use contact_19  contact_19_122
timestamp 1634918361
transform 1 0 1726 0 1 19200
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1634918361
transform 1 0 1729 0 1 19199
box 0 0 1 1
use contact_13  contact_13_122
timestamp 1634918361
transform 1 0 1733 0 1 19191
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1634918361
transform 1 0 1725 0 1 18859
box 0 0 1 1
use contact_19  contact_19_123
timestamp 1634918361
transform 1 0 1726 0 1 18864
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1634918361
transform 1 0 1729 0 1 18863
box 0 0 1 1
use contact_13  contact_13_123
timestamp 1634918361
transform 1 0 1733 0 1 18855
box 0 0 1 1
use contact_19  contact_19_124
timestamp 1634918361
transform 1 0 1726 0 1 18528
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1634918361
transform 1 0 1729 0 1 18527
box 0 0 1 1
use contact_13  contact_13_124
timestamp 1634918361
transform 1 0 1733 0 1 18519
box 0 0 1 1
use contact_19  contact_19_125
timestamp 1634918361
transform 1 0 1726 0 1 18192
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1634918361
transform 1 0 1729 0 1 18191
box 0 0 1 1
use contact_13  contact_13_125
timestamp 1634918361
transform 1 0 1733 0 1 18183
box 0 0 1 1
use contact_19  contact_19_126
timestamp 1634918361
transform 1 0 1726 0 1 17856
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1634918361
transform 1 0 1729 0 1 17855
box 0 0 1 1
use contact_13  contact_13_126
timestamp 1634918361
transform 1 0 1733 0 1 17847
box 0 0 1 1
use contact_19  contact_19_127
timestamp 1634918361
transform 1 0 1726 0 1 17520
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1634918361
transform 1 0 1729 0 1 17519
box 0 0 1 1
use contact_13  contact_13_127
timestamp 1634918361
transform 1 0 1733 0 1 17511
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1634918361
transform 1 0 1725 0 1 17179
box 0 0 1 1
use contact_19  contact_19_128
timestamp 1634918361
transform 1 0 1726 0 1 17184
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1634918361
transform 1 0 1729 0 1 17183
box 0 0 1 1
use contact_13  contact_13_128
timestamp 1634918361
transform 1 0 1733 0 1 17175
box 0 0 1 1
use contact_19  contact_19_129
timestamp 1634918361
transform 1 0 1726 0 1 16848
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1634918361
transform 1 0 1729 0 1 16847
box 0 0 1 1
use contact_13  contact_13_129
timestamp 1634918361
transform 1 0 1733 0 1 16839
box 0 0 1 1
use contact_19  contact_19_130
timestamp 1634918361
transform 1 0 1726 0 1 16512
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1634918361
transform 1 0 1729 0 1 16511
box 0 0 1 1
use contact_13  contact_13_130
timestamp 1634918361
transform 1 0 1733 0 1 16503
box 0 0 1 1
use contact_19  contact_19_131
timestamp 1634918361
transform 1 0 1726 0 1 16176
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1634918361
transform 1 0 1729 0 1 16175
box 0 0 1 1
use contact_13  contact_13_131
timestamp 1634918361
transform 1 0 1733 0 1 16167
box 0 0 1 1
use contact_19  contact_19_132
timestamp 1634918361
transform 1 0 1726 0 1 15840
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1634918361
transform 1 0 1729 0 1 15839
box 0 0 1 1
use contact_13  contact_13_132
timestamp 1634918361
transform 1 0 1733 0 1 15831
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1634918361
transform 1 0 1725 0 1 15499
box 0 0 1 1
use contact_19  contact_19_133
timestamp 1634918361
transform 1 0 1726 0 1 15504
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1634918361
transform 1 0 1729 0 1 15503
box 0 0 1 1
use contact_13  contact_13_133
timestamp 1634918361
transform 1 0 1733 0 1 15495
box 0 0 1 1
use contact_19  contact_19_134
timestamp 1634918361
transform 1 0 1726 0 1 15168
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1634918361
transform 1 0 1729 0 1 15167
box 0 0 1 1
use contact_13  contact_13_134
timestamp 1634918361
transform 1 0 1733 0 1 15159
box 0 0 1 1
use contact_19  contact_19_135
timestamp 1634918361
transform 1 0 1726 0 1 14832
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1634918361
transform 1 0 1729 0 1 14831
box 0 0 1 1
use contact_13  contact_13_135
timestamp 1634918361
transform 1 0 1733 0 1 14823
box 0 0 1 1
use contact_19  contact_19_136
timestamp 1634918361
transform 1 0 1726 0 1 14496
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1634918361
transform 1 0 1729 0 1 14495
box 0 0 1 1
use contact_13  contact_13_136
timestamp 1634918361
transform 1 0 1733 0 1 14487
box 0 0 1 1
use contact_19  contact_19_137
timestamp 1634918361
transform 1 0 1726 0 1 14160
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1634918361
transform 1 0 1729 0 1 14159
box 0 0 1 1
use contact_13  contact_13_137
timestamp 1634918361
transform 1 0 1733 0 1 14151
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1634918361
transform 1 0 1725 0 1 13819
box 0 0 1 1
use contact_19  contact_19_138
timestamp 1634918361
transform 1 0 1726 0 1 13824
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1634918361
transform 1 0 1729 0 1 13823
box 0 0 1 1
use contact_13  contact_13_138
timestamp 1634918361
transform 1 0 1733 0 1 13815
box 0 0 1 1
use contact_19  contact_19_139
timestamp 1634918361
transform 1 0 1726 0 1 13488
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1634918361
transform 1 0 1729 0 1 13487
box 0 0 1 1
use contact_13  contact_13_139
timestamp 1634918361
transform 1 0 1733 0 1 13479
box 0 0 1 1
use contact_19  contact_19_140
timestamp 1634918361
transform 1 0 1726 0 1 13152
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1634918361
transform 1 0 1729 0 1 13151
box 0 0 1 1
use contact_13  contact_13_140
timestamp 1634918361
transform 1 0 1733 0 1 13143
box 0 0 1 1
use contact_19  contact_19_141
timestamp 1634918361
transform 1 0 1726 0 1 12816
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1634918361
transform 1 0 1729 0 1 12815
box 0 0 1 1
use contact_13  contact_13_141
timestamp 1634918361
transform 1 0 1733 0 1 12807
box 0 0 1 1
use contact_19  contact_19_142
timestamp 1634918361
transform 1 0 1726 0 1 12480
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1634918361
transform 1 0 1729 0 1 12479
box 0 0 1 1
use contact_13  contact_13_142
timestamp 1634918361
transform 1 0 1733 0 1 12471
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1634918361
transform 1 0 1725 0 1 12139
box 0 0 1 1
use contact_19  contact_19_143
timestamp 1634918361
transform 1 0 1726 0 1 12144
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1634918361
transform 1 0 1729 0 1 12143
box 0 0 1 1
use contact_13  contact_13_143
timestamp 1634918361
transform 1 0 1733 0 1 12135
box 0 0 1 1
use contact_19  contact_19_144
timestamp 1634918361
transform 1 0 1726 0 1 11808
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1634918361
transform 1 0 1729 0 1 11807
box 0 0 1 1
use contact_13  contact_13_144
timestamp 1634918361
transform 1 0 1733 0 1 11799
box 0 0 1 1
use contact_19  contact_19_145
timestamp 1634918361
transform 1 0 1726 0 1 11472
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1634918361
transform 1 0 1729 0 1 11471
box 0 0 1 1
use contact_13  contact_13_145
timestamp 1634918361
transform 1 0 1733 0 1 11463
box 0 0 1 1
use contact_19  contact_19_146
timestamp 1634918361
transform 1 0 1726 0 1 11136
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1634918361
transform 1 0 1729 0 1 11135
box 0 0 1 1
use contact_13  contact_13_146
timestamp 1634918361
transform 1 0 1733 0 1 11127
box 0 0 1 1
use contact_19  contact_19_147
timestamp 1634918361
transform 1 0 1726 0 1 10800
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1634918361
transform 1 0 1729 0 1 10799
box 0 0 1 1
use contact_13  contact_13_147
timestamp 1634918361
transform 1 0 1733 0 1 10791
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1634918361
transform 1 0 1725 0 1 10459
box 0 0 1 1
use contact_19  contact_19_148
timestamp 1634918361
transform 1 0 1726 0 1 10464
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1634918361
transform 1 0 1729 0 1 10463
box 0 0 1 1
use contact_13  contact_13_148
timestamp 1634918361
transform 1 0 1733 0 1 10455
box 0 0 1 1
use contact_19  contact_19_149
timestamp 1634918361
transform 1 0 1726 0 1 10128
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1634918361
transform 1 0 1729 0 1 10127
box 0 0 1 1
use contact_13  contact_13_149
timestamp 1634918361
transform 1 0 1733 0 1 10119
box 0 0 1 1
use contact_19  contact_19_150
timestamp 1634918361
transform 1 0 1726 0 1 9792
box 0 0 1 1
use contact_14  contact_14_150
timestamp 1634918361
transform 1 0 1729 0 1 9791
box 0 0 1 1
use contact_13  contact_13_150
timestamp 1634918361
transform 1 0 1733 0 1 9783
box 0 0 1 1
use contact_19  contact_19_151
timestamp 1634918361
transform 1 0 1726 0 1 9456
box 0 0 1 1
use contact_14  contact_14_151
timestamp 1634918361
transform 1 0 1729 0 1 9455
box 0 0 1 1
use contact_13  contact_13_151
timestamp 1634918361
transform 1 0 1733 0 1 9447
box 0 0 1 1
use contact_19  contact_19_152
timestamp 1634918361
transform 1 0 1726 0 1 9120
box 0 0 1 1
use contact_14  contact_14_152
timestamp 1634918361
transform 1 0 1729 0 1 9119
box 0 0 1 1
use contact_13  contact_13_152
timestamp 1634918361
transform 1 0 1733 0 1 9111
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1634918361
transform 1 0 1725 0 1 8779
box 0 0 1 1
use contact_19  contact_19_153
timestamp 1634918361
transform 1 0 1726 0 1 8784
box 0 0 1 1
use contact_14  contact_14_153
timestamp 1634918361
transform 1 0 1729 0 1 8783
box 0 0 1 1
use contact_13  contact_13_153
timestamp 1634918361
transform 1 0 1733 0 1 8775
box 0 0 1 1
use contact_19  contact_19_154
timestamp 1634918361
transform 1 0 1726 0 1 8448
box 0 0 1 1
use contact_14  contact_14_154
timestamp 1634918361
transform 1 0 1729 0 1 8447
box 0 0 1 1
use contact_13  contact_13_154
timestamp 1634918361
transform 1 0 1733 0 1 8439
box 0 0 1 1
use contact_19  contact_19_155
timestamp 1634918361
transform 1 0 1726 0 1 8112
box 0 0 1 1
use contact_14  contact_14_155
timestamp 1634918361
transform 1 0 1729 0 1 8111
box 0 0 1 1
use contact_13  contact_13_155
timestamp 1634918361
transform 1 0 1733 0 1 8103
box 0 0 1 1
use contact_19  contact_19_156
timestamp 1634918361
transform 1 0 1726 0 1 7776
box 0 0 1 1
use contact_14  contact_14_156
timestamp 1634918361
transform 1 0 1729 0 1 7775
box 0 0 1 1
use contact_13  contact_13_156
timestamp 1634918361
transform 1 0 1733 0 1 7767
box 0 0 1 1
use contact_19  contact_19_157
timestamp 1634918361
transform 1 0 1726 0 1 7440
box 0 0 1 1
use contact_14  contact_14_157
timestamp 1634918361
transform 1 0 1729 0 1 7439
box 0 0 1 1
use contact_13  contact_13_157
timestamp 1634918361
transform 1 0 1733 0 1 7431
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1634918361
transform 1 0 1725 0 1 7099
box 0 0 1 1
use contact_19  contact_19_158
timestamp 1634918361
transform 1 0 1726 0 1 7104
box 0 0 1 1
use contact_14  contact_14_158
timestamp 1634918361
transform 1 0 1729 0 1 7103
box 0 0 1 1
use contact_13  contact_13_158
timestamp 1634918361
transform 1 0 1733 0 1 7095
box 0 0 1 1
use contact_19  contact_19_159
timestamp 1634918361
transform 1 0 1726 0 1 6768
box 0 0 1 1
use contact_14  contact_14_159
timestamp 1634918361
transform 1 0 1729 0 1 6767
box 0 0 1 1
use contact_13  contact_13_159
timestamp 1634918361
transform 1 0 1733 0 1 6759
box 0 0 1 1
use contact_19  contact_19_160
timestamp 1634918361
transform 1 0 1726 0 1 6432
box 0 0 1 1
use contact_14  contact_14_160
timestamp 1634918361
transform 1 0 1729 0 1 6431
box 0 0 1 1
use contact_13  contact_13_160
timestamp 1634918361
transform 1 0 1733 0 1 6423
box 0 0 1 1
use contact_19  contact_19_161
timestamp 1634918361
transform 1 0 1726 0 1 6096
box 0 0 1 1
use contact_14  contact_14_161
timestamp 1634918361
transform 1 0 1729 0 1 6095
box 0 0 1 1
use contact_13  contact_13_161
timestamp 1634918361
transform 1 0 1733 0 1 6087
box 0 0 1 1
use contact_19  contact_19_162
timestamp 1634918361
transform 1 0 1726 0 1 5760
box 0 0 1 1
use contact_14  contact_14_162
timestamp 1634918361
transform 1 0 1729 0 1 5759
box 0 0 1 1
use contact_13  contact_13_162
timestamp 1634918361
transform 1 0 1733 0 1 5751
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1634918361
transform 1 0 1725 0 1 5419
box 0 0 1 1
use contact_19  contact_19_163
timestamp 1634918361
transform 1 0 1726 0 1 5424
box 0 0 1 1
use contact_14  contact_14_163
timestamp 1634918361
transform 1 0 1729 0 1 5423
box 0 0 1 1
use contact_13  contact_13_163
timestamp 1634918361
transform 1 0 1733 0 1 5415
box 0 0 1 1
use contact_19  contact_19_164
timestamp 1634918361
transform 1 0 1726 0 1 5088
box 0 0 1 1
use contact_14  contact_14_164
timestamp 1634918361
transform 1 0 1729 0 1 5087
box 0 0 1 1
use contact_13  contact_13_164
timestamp 1634918361
transform 1 0 1733 0 1 5079
box 0 0 1 1
use contact_19  contact_19_165
timestamp 1634918361
transform 1 0 1726 0 1 4752
box 0 0 1 1
use contact_14  contact_14_165
timestamp 1634918361
transform 1 0 1729 0 1 4751
box 0 0 1 1
use contact_13  contact_13_165
timestamp 1634918361
transform 1 0 1733 0 1 4743
box 0 0 1 1
use contact_19  contact_19_166
timestamp 1634918361
transform 1 0 1726 0 1 4416
box 0 0 1 1
use contact_14  contact_14_166
timestamp 1634918361
transform 1 0 1729 0 1 4415
box 0 0 1 1
use contact_13  contact_13_166
timestamp 1634918361
transform 1 0 1733 0 1 4407
box 0 0 1 1
use contact_19  contact_19_167
timestamp 1634918361
transform 1 0 1726 0 1 4080
box 0 0 1 1
use contact_14  contact_14_167
timestamp 1634918361
transform 1 0 1729 0 1 4079
box 0 0 1 1
use contact_13  contact_13_167
timestamp 1634918361
transform 1 0 1733 0 1 4071
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1634918361
transform 1 0 1725 0 1 3739
box 0 0 1 1
use contact_19  contact_19_168
timestamp 1634918361
transform 1 0 1726 0 1 3744
box 0 0 1 1
use contact_14  contact_14_168
timestamp 1634918361
transform 1 0 1729 0 1 3743
box 0 0 1 1
use contact_13  contact_13_168
timestamp 1634918361
transform 1 0 1733 0 1 3735
box 0 0 1 1
use contact_19  contact_19_169
timestamp 1634918361
transform 1 0 1726 0 1 3408
box 0 0 1 1
use contact_14  contact_14_169
timestamp 1634918361
transform 1 0 1729 0 1 3407
box 0 0 1 1
use contact_13  contact_13_169
timestamp 1634918361
transform 1 0 1733 0 1 3399
box 0 0 1 1
use contact_19  contact_19_170
timestamp 1634918361
transform 1 0 1726 0 1 3072
box 0 0 1 1
use contact_14  contact_14_170
timestamp 1634918361
transform 1 0 1729 0 1 3071
box 0 0 1 1
use contact_13  contact_13_170
timestamp 1634918361
transform 1 0 1733 0 1 3063
box 0 0 1 1
use contact_19  contact_19_171
timestamp 1634918361
transform 1 0 1726 0 1 2736
box 0 0 1 1
use contact_14  contact_14_171
timestamp 1634918361
transform 1 0 1729 0 1 2735
box 0 0 1 1
use contact_13  contact_13_171
timestamp 1634918361
transform 1 0 1733 0 1 2727
box 0 0 1 1
use contact_19  contact_19_172
timestamp 1634918361
transform 1 0 1726 0 1 2400
box 0 0 1 1
use contact_14  contact_14_172
timestamp 1634918361
transform 1 0 1729 0 1 2399
box 0 0 1 1
use contact_13  contact_13_172
timestamp 1634918361
transform 1 0 1733 0 1 2391
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1634918361
transform 1 0 1725 0 1 2059
box 0 0 1 1
use contact_19  contact_19_173
timestamp 1634918361
transform 1 0 1726 0 1 2064
box 0 0 1 1
use contact_14  contact_14_173
timestamp 1634918361
transform 1 0 1729 0 1 2063
box 0 0 1 1
use contact_13  contact_13_173
timestamp 1634918361
transform 1 0 1733 0 1 2055
box 0 0 1 1
use contact_14  contact_14_174
timestamp 1634918361
transform 1 0 41041 0 1 31351
box 0 0 1 1
use contact_13  contact_13_174
timestamp 1634918361
transform 1 0 41045 0 1 31343
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1634918361
transform 1 0 40701 0 1 31347
box 0 0 1 1
use contact_19  contact_19_174
timestamp 1634918361
transform 1 0 40702 0 1 31352
box 0 0 1 1
use contact_14  contact_14_175
timestamp 1634918361
transform 1 0 40705 0 1 31351
box 0 0 1 1
use contact_13  contact_13_175
timestamp 1634918361
transform 1 0 40709 0 1 31343
box 0 0 1 1
use contact_14  contact_14_176
timestamp 1634918361
transform 1 0 40369 0 1 31351
box 0 0 1 1
use contact_13  contact_13_176
timestamp 1634918361
transform 1 0 40373 0 1 31343
box 0 0 1 1
use contact_14  contact_14_177
timestamp 1634918361
transform 1 0 40033 0 1 31351
box 0 0 1 1
use contact_13  contact_13_177
timestamp 1634918361
transform 1 0 40037 0 1 31343
box 0 0 1 1
use contact_14  contact_14_178
timestamp 1634918361
transform 1 0 39697 0 1 31351
box 0 0 1 1
use contact_13  contact_13_178
timestamp 1634918361
transform 1 0 39701 0 1 31343
box 0 0 1 1
use contact_14  contact_14_179
timestamp 1634918361
transform 1 0 39361 0 1 31351
box 0 0 1 1
use contact_13  contact_13_179
timestamp 1634918361
transform 1 0 39365 0 1 31343
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1634918361
transform 1 0 39021 0 1 31347
box 0 0 1 1
use contact_19  contact_19_175
timestamp 1634918361
transform 1 0 39022 0 1 31352
box 0 0 1 1
use contact_14  contact_14_180
timestamp 1634918361
transform 1 0 39025 0 1 31351
box 0 0 1 1
use contact_13  contact_13_180
timestamp 1634918361
transform 1 0 39029 0 1 31343
box 0 0 1 1
use contact_14  contact_14_181
timestamp 1634918361
transform 1 0 38689 0 1 31351
box 0 0 1 1
use contact_13  contact_13_181
timestamp 1634918361
transform 1 0 38693 0 1 31343
box 0 0 1 1
use contact_14  contact_14_182
timestamp 1634918361
transform 1 0 38353 0 1 31351
box 0 0 1 1
use contact_13  contact_13_182
timestamp 1634918361
transform 1 0 38357 0 1 31343
box 0 0 1 1
use contact_14  contact_14_183
timestamp 1634918361
transform 1 0 38017 0 1 31351
box 0 0 1 1
use contact_13  contact_13_183
timestamp 1634918361
transform 1 0 38021 0 1 31343
box 0 0 1 1
use contact_14  contact_14_184
timestamp 1634918361
transform 1 0 37681 0 1 31351
box 0 0 1 1
use contact_13  contact_13_184
timestamp 1634918361
transform 1 0 37685 0 1 31343
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1634918361
transform 1 0 37341 0 1 31347
box 0 0 1 1
use contact_19  contact_19_176
timestamp 1634918361
transform 1 0 37342 0 1 31352
box 0 0 1 1
use contact_14  contact_14_185
timestamp 1634918361
transform 1 0 37345 0 1 31351
box 0 0 1 1
use contact_13  contact_13_185
timestamp 1634918361
transform 1 0 37349 0 1 31343
box 0 0 1 1
use contact_14  contact_14_186
timestamp 1634918361
transform 1 0 37009 0 1 31351
box 0 0 1 1
use contact_13  contact_13_186
timestamp 1634918361
transform 1 0 37013 0 1 31343
box 0 0 1 1
use contact_14  contact_14_187
timestamp 1634918361
transform 1 0 36673 0 1 31351
box 0 0 1 1
use contact_13  contact_13_187
timestamp 1634918361
transform 1 0 36677 0 1 31343
box 0 0 1 1
use contact_14  contact_14_188
timestamp 1634918361
transform 1 0 36337 0 1 31351
box 0 0 1 1
use contact_13  contact_13_188
timestamp 1634918361
transform 1 0 36341 0 1 31343
box 0 0 1 1
use contact_14  contact_14_189
timestamp 1634918361
transform 1 0 36001 0 1 31351
box 0 0 1 1
use contact_13  contact_13_189
timestamp 1634918361
transform 1 0 36005 0 1 31343
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1634918361
transform 1 0 35661 0 1 31347
box 0 0 1 1
use contact_19  contact_19_177
timestamp 1634918361
transform 1 0 35662 0 1 31352
box 0 0 1 1
use contact_14  contact_14_190
timestamp 1634918361
transform 1 0 35665 0 1 31351
box 0 0 1 1
use contact_13  contact_13_190
timestamp 1634918361
transform 1 0 35669 0 1 31343
box 0 0 1 1
use contact_14  contact_14_191
timestamp 1634918361
transform 1 0 35329 0 1 31351
box 0 0 1 1
use contact_13  contact_13_191
timestamp 1634918361
transform 1 0 35333 0 1 31343
box 0 0 1 1
use contact_14  contact_14_192
timestamp 1634918361
transform 1 0 34993 0 1 31351
box 0 0 1 1
use contact_13  contact_13_192
timestamp 1634918361
transform 1 0 34997 0 1 31343
box 0 0 1 1
use contact_14  contact_14_193
timestamp 1634918361
transform 1 0 34657 0 1 31351
box 0 0 1 1
use contact_13  contact_13_193
timestamp 1634918361
transform 1 0 34661 0 1 31343
box 0 0 1 1
use contact_14  contact_14_194
timestamp 1634918361
transform 1 0 34321 0 1 31351
box 0 0 1 1
use contact_13  contact_13_194
timestamp 1634918361
transform 1 0 34325 0 1 31343
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1634918361
transform 1 0 33981 0 1 31347
box 0 0 1 1
use contact_19  contact_19_178
timestamp 1634918361
transform 1 0 33982 0 1 31352
box 0 0 1 1
use contact_14  contact_14_195
timestamp 1634918361
transform 1 0 33985 0 1 31351
box 0 0 1 1
use contact_13  contact_13_195
timestamp 1634918361
transform 1 0 33989 0 1 31343
box 0 0 1 1
use contact_14  contact_14_196
timestamp 1634918361
transform 1 0 33649 0 1 31351
box 0 0 1 1
use contact_13  contact_13_196
timestamp 1634918361
transform 1 0 33653 0 1 31343
box 0 0 1 1
use contact_14  contact_14_197
timestamp 1634918361
transform 1 0 33313 0 1 31351
box 0 0 1 1
use contact_13  contact_13_197
timestamp 1634918361
transform 1 0 33317 0 1 31343
box 0 0 1 1
use contact_14  contact_14_198
timestamp 1634918361
transform 1 0 32977 0 1 31351
box 0 0 1 1
use contact_13  contact_13_198
timestamp 1634918361
transform 1 0 32981 0 1 31343
box 0 0 1 1
use contact_14  contact_14_199
timestamp 1634918361
transform 1 0 32641 0 1 31351
box 0 0 1 1
use contact_13  contact_13_199
timestamp 1634918361
transform 1 0 32645 0 1 31343
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1634918361
transform 1 0 32301 0 1 31347
box 0 0 1 1
use contact_19  contact_19_179
timestamp 1634918361
transform 1 0 32302 0 1 31352
box 0 0 1 1
use contact_14  contact_14_200
timestamp 1634918361
transform 1 0 32305 0 1 31351
box 0 0 1 1
use contact_13  contact_13_200
timestamp 1634918361
transform 1 0 32309 0 1 31343
box 0 0 1 1
use contact_14  contact_14_201
timestamp 1634918361
transform 1 0 31969 0 1 31351
box 0 0 1 1
use contact_13  contact_13_201
timestamp 1634918361
transform 1 0 31973 0 1 31343
box 0 0 1 1
use contact_14  contact_14_202
timestamp 1634918361
transform 1 0 31633 0 1 31351
box 0 0 1 1
use contact_13  contact_13_202
timestamp 1634918361
transform 1 0 31637 0 1 31343
box 0 0 1 1
use contact_14  contact_14_203
timestamp 1634918361
transform 1 0 31297 0 1 31351
box 0 0 1 1
use contact_13  contact_13_203
timestamp 1634918361
transform 1 0 31301 0 1 31343
box 0 0 1 1
use contact_14  contact_14_204
timestamp 1634918361
transform 1 0 30961 0 1 31351
box 0 0 1 1
use contact_13  contact_13_204
timestamp 1634918361
transform 1 0 30965 0 1 31343
box 0 0 1 1
use contact_7  contact_7_42
timestamp 1634918361
transform 1 0 30621 0 1 31347
box 0 0 1 1
use contact_19  contact_19_180
timestamp 1634918361
transform 1 0 30622 0 1 31352
box 0 0 1 1
use contact_14  contact_14_205
timestamp 1634918361
transform 1 0 30625 0 1 31351
box 0 0 1 1
use contact_13  contact_13_205
timestamp 1634918361
transform 1 0 30629 0 1 31343
box 0 0 1 1
use contact_14  contact_14_206
timestamp 1634918361
transform 1 0 30289 0 1 31351
box 0 0 1 1
use contact_13  contact_13_206
timestamp 1634918361
transform 1 0 30293 0 1 31343
box 0 0 1 1
use contact_14  contact_14_207
timestamp 1634918361
transform 1 0 29953 0 1 31351
box 0 0 1 1
use contact_13  contact_13_207
timestamp 1634918361
transform 1 0 29957 0 1 31343
box 0 0 1 1
use contact_14  contact_14_208
timestamp 1634918361
transform 1 0 29617 0 1 31351
box 0 0 1 1
use contact_13  contact_13_208
timestamp 1634918361
transform 1 0 29621 0 1 31343
box 0 0 1 1
use contact_14  contact_14_209
timestamp 1634918361
transform 1 0 29281 0 1 31351
box 0 0 1 1
use contact_13  contact_13_209
timestamp 1634918361
transform 1 0 29285 0 1 31343
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1634918361
transform 1 0 28941 0 1 31347
box 0 0 1 1
use contact_19  contact_19_181
timestamp 1634918361
transform 1 0 28942 0 1 31352
box 0 0 1 1
use contact_14  contact_14_210
timestamp 1634918361
transform 1 0 28945 0 1 31351
box 0 0 1 1
use contact_13  contact_13_210
timestamp 1634918361
transform 1 0 28949 0 1 31343
box 0 0 1 1
use contact_14  contact_14_211
timestamp 1634918361
transform 1 0 28609 0 1 31351
box 0 0 1 1
use contact_13  contact_13_211
timestamp 1634918361
transform 1 0 28613 0 1 31343
box 0 0 1 1
use contact_14  contact_14_212
timestamp 1634918361
transform 1 0 28273 0 1 31351
box 0 0 1 1
use contact_13  contact_13_212
timestamp 1634918361
transform 1 0 28277 0 1 31343
box 0 0 1 1
use contact_14  contact_14_213
timestamp 1634918361
transform 1 0 27937 0 1 31351
box 0 0 1 1
use contact_13  contact_13_213
timestamp 1634918361
transform 1 0 27941 0 1 31343
box 0 0 1 1
use contact_14  contact_14_214
timestamp 1634918361
transform 1 0 27601 0 1 31351
box 0 0 1 1
use contact_13  contact_13_214
timestamp 1634918361
transform 1 0 27605 0 1 31343
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1634918361
transform 1 0 27261 0 1 31347
box 0 0 1 1
use contact_19  contact_19_182
timestamp 1634918361
transform 1 0 27262 0 1 31352
box 0 0 1 1
use contact_14  contact_14_215
timestamp 1634918361
transform 1 0 27265 0 1 31351
box 0 0 1 1
use contact_13  contact_13_215
timestamp 1634918361
transform 1 0 27269 0 1 31343
box 0 0 1 1
use contact_14  contact_14_216
timestamp 1634918361
transform 1 0 26929 0 1 31351
box 0 0 1 1
use contact_13  contact_13_216
timestamp 1634918361
transform 1 0 26933 0 1 31343
box 0 0 1 1
use contact_14  contact_14_217
timestamp 1634918361
transform 1 0 26593 0 1 31351
box 0 0 1 1
use contact_13  contact_13_217
timestamp 1634918361
transform 1 0 26597 0 1 31343
box 0 0 1 1
use contact_14  contact_14_218
timestamp 1634918361
transform 1 0 26257 0 1 31351
box 0 0 1 1
use contact_13  contact_13_218
timestamp 1634918361
transform 1 0 26261 0 1 31343
box 0 0 1 1
use contact_14  contact_14_219
timestamp 1634918361
transform 1 0 25921 0 1 31351
box 0 0 1 1
use contact_13  contact_13_219
timestamp 1634918361
transform 1 0 25925 0 1 31343
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1634918361
transform 1 0 25581 0 1 31347
box 0 0 1 1
use contact_19  contact_19_183
timestamp 1634918361
transform 1 0 25582 0 1 31352
box 0 0 1 1
use contact_14  contact_14_220
timestamp 1634918361
transform 1 0 25585 0 1 31351
box 0 0 1 1
use contact_13  contact_13_220
timestamp 1634918361
transform 1 0 25589 0 1 31343
box 0 0 1 1
use contact_14  contact_14_221
timestamp 1634918361
transform 1 0 25249 0 1 31351
box 0 0 1 1
use contact_13  contact_13_221
timestamp 1634918361
transform 1 0 25253 0 1 31343
box 0 0 1 1
use contact_14  contact_14_222
timestamp 1634918361
transform 1 0 24913 0 1 31351
box 0 0 1 1
use contact_13  contact_13_222
timestamp 1634918361
transform 1 0 24917 0 1 31343
box 0 0 1 1
use contact_14  contact_14_223
timestamp 1634918361
transform 1 0 24577 0 1 31351
box 0 0 1 1
use contact_13  contact_13_223
timestamp 1634918361
transform 1 0 24581 0 1 31343
box 0 0 1 1
use contact_14  contact_14_224
timestamp 1634918361
transform 1 0 24241 0 1 31351
box 0 0 1 1
use contact_13  contact_13_224
timestamp 1634918361
transform 1 0 24245 0 1 31343
box 0 0 1 1
use contact_7  contact_7_46
timestamp 1634918361
transform 1 0 23901 0 1 31347
box 0 0 1 1
use contact_19  contact_19_184
timestamp 1634918361
transform 1 0 23902 0 1 31352
box 0 0 1 1
use contact_14  contact_14_225
timestamp 1634918361
transform 1 0 23905 0 1 31351
box 0 0 1 1
use contact_13  contact_13_225
timestamp 1634918361
transform 1 0 23909 0 1 31343
box 0 0 1 1
use contact_14  contact_14_226
timestamp 1634918361
transform 1 0 23569 0 1 31351
box 0 0 1 1
use contact_13  contact_13_226
timestamp 1634918361
transform 1 0 23573 0 1 31343
box 0 0 1 1
use contact_14  contact_14_227
timestamp 1634918361
transform 1 0 23233 0 1 31351
box 0 0 1 1
use contact_13  contact_13_227
timestamp 1634918361
transform 1 0 23237 0 1 31343
box 0 0 1 1
use contact_14  contact_14_228
timestamp 1634918361
transform 1 0 22897 0 1 31351
box 0 0 1 1
use contact_13  contact_13_228
timestamp 1634918361
transform 1 0 22901 0 1 31343
box 0 0 1 1
use contact_14  contact_14_229
timestamp 1634918361
transform 1 0 22561 0 1 31351
box 0 0 1 1
use contact_13  contact_13_229
timestamp 1634918361
transform 1 0 22565 0 1 31343
box 0 0 1 1
use contact_7  contact_7_47
timestamp 1634918361
transform 1 0 22221 0 1 31347
box 0 0 1 1
use contact_19  contact_19_185
timestamp 1634918361
transform 1 0 22222 0 1 31352
box 0 0 1 1
use contact_14  contact_14_230
timestamp 1634918361
transform 1 0 22225 0 1 31351
box 0 0 1 1
use contact_13  contact_13_230
timestamp 1634918361
transform 1 0 22229 0 1 31343
box 0 0 1 1
use contact_14  contact_14_231
timestamp 1634918361
transform 1 0 21889 0 1 31351
box 0 0 1 1
use contact_13  contact_13_231
timestamp 1634918361
transform 1 0 21893 0 1 31343
box 0 0 1 1
use contact_14  contact_14_232
timestamp 1634918361
transform 1 0 21553 0 1 31351
box 0 0 1 1
use contact_13  contact_13_232
timestamp 1634918361
transform 1 0 21557 0 1 31343
box 0 0 1 1
use contact_14  contact_14_233
timestamp 1634918361
transform 1 0 21217 0 1 31351
box 0 0 1 1
use contact_13  contact_13_233
timestamp 1634918361
transform 1 0 21221 0 1 31343
box 0 0 1 1
use contact_14  contact_14_234
timestamp 1634918361
transform 1 0 20881 0 1 31351
box 0 0 1 1
use contact_13  contact_13_234
timestamp 1634918361
transform 1 0 20885 0 1 31343
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1634918361
transform 1 0 20541 0 1 31347
box 0 0 1 1
use contact_19  contact_19_186
timestamp 1634918361
transform 1 0 20542 0 1 31352
box 0 0 1 1
use contact_14  contact_14_235
timestamp 1634918361
transform 1 0 20545 0 1 31351
box 0 0 1 1
use contact_13  contact_13_235
timestamp 1634918361
transform 1 0 20549 0 1 31343
box 0 0 1 1
use contact_14  contact_14_236
timestamp 1634918361
transform 1 0 20209 0 1 31351
box 0 0 1 1
use contact_13  contact_13_236
timestamp 1634918361
transform 1 0 20213 0 1 31343
box 0 0 1 1
use contact_14  contact_14_237
timestamp 1634918361
transform 1 0 19873 0 1 31351
box 0 0 1 1
use contact_13  contact_13_237
timestamp 1634918361
transform 1 0 19877 0 1 31343
box 0 0 1 1
use contact_14  contact_14_238
timestamp 1634918361
transform 1 0 19537 0 1 31351
box 0 0 1 1
use contact_13  contact_13_238
timestamp 1634918361
transform 1 0 19541 0 1 31343
box 0 0 1 1
use contact_14  contact_14_239
timestamp 1634918361
transform 1 0 19201 0 1 31351
box 0 0 1 1
use contact_13  contact_13_239
timestamp 1634918361
transform 1 0 19205 0 1 31343
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1634918361
transform 1 0 18861 0 1 31347
box 0 0 1 1
use contact_19  contact_19_187
timestamp 1634918361
transform 1 0 18862 0 1 31352
box 0 0 1 1
use contact_14  contact_14_240
timestamp 1634918361
transform 1 0 18865 0 1 31351
box 0 0 1 1
use contact_13  contact_13_240
timestamp 1634918361
transform 1 0 18869 0 1 31343
box 0 0 1 1
use contact_14  contact_14_241
timestamp 1634918361
transform 1 0 18529 0 1 31351
box 0 0 1 1
use contact_13  contact_13_241
timestamp 1634918361
transform 1 0 18533 0 1 31343
box 0 0 1 1
use contact_14  contact_14_242
timestamp 1634918361
transform 1 0 18193 0 1 31351
box 0 0 1 1
use contact_13  contact_13_242
timestamp 1634918361
transform 1 0 18197 0 1 31343
box 0 0 1 1
use contact_14  contact_14_243
timestamp 1634918361
transform 1 0 17857 0 1 31351
box 0 0 1 1
use contact_13  contact_13_243
timestamp 1634918361
transform 1 0 17861 0 1 31343
box 0 0 1 1
use contact_14  contact_14_244
timestamp 1634918361
transform 1 0 17521 0 1 31351
box 0 0 1 1
use contact_13  contact_13_244
timestamp 1634918361
transform 1 0 17525 0 1 31343
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1634918361
transform 1 0 17181 0 1 31347
box 0 0 1 1
use contact_19  contact_19_188
timestamp 1634918361
transform 1 0 17182 0 1 31352
box 0 0 1 1
use contact_14  contact_14_245
timestamp 1634918361
transform 1 0 17185 0 1 31351
box 0 0 1 1
use contact_13  contact_13_245
timestamp 1634918361
transform 1 0 17189 0 1 31343
box 0 0 1 1
use contact_14  contact_14_246
timestamp 1634918361
transform 1 0 16849 0 1 31351
box 0 0 1 1
use contact_13  contact_13_246
timestamp 1634918361
transform 1 0 16853 0 1 31343
box 0 0 1 1
use contact_14  contact_14_247
timestamp 1634918361
transform 1 0 16513 0 1 31351
box 0 0 1 1
use contact_13  contact_13_247
timestamp 1634918361
transform 1 0 16517 0 1 31343
box 0 0 1 1
use contact_14  contact_14_248
timestamp 1634918361
transform 1 0 16177 0 1 31351
box 0 0 1 1
use contact_13  contact_13_248
timestamp 1634918361
transform 1 0 16181 0 1 31343
box 0 0 1 1
use contact_14  contact_14_249
timestamp 1634918361
transform 1 0 15841 0 1 31351
box 0 0 1 1
use contact_13  contact_13_249
timestamp 1634918361
transform 1 0 15845 0 1 31343
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1634918361
transform 1 0 15501 0 1 31347
box 0 0 1 1
use contact_19  contact_19_189
timestamp 1634918361
transform 1 0 15502 0 1 31352
box 0 0 1 1
use contact_14  contact_14_250
timestamp 1634918361
transform 1 0 15505 0 1 31351
box 0 0 1 1
use contact_13  contact_13_250
timestamp 1634918361
transform 1 0 15509 0 1 31343
box 0 0 1 1
use contact_14  contact_14_251
timestamp 1634918361
transform 1 0 15169 0 1 31351
box 0 0 1 1
use contact_13  contact_13_251
timestamp 1634918361
transform 1 0 15173 0 1 31343
box 0 0 1 1
use contact_14  contact_14_252
timestamp 1634918361
transform 1 0 14833 0 1 31351
box 0 0 1 1
use contact_13  contact_13_252
timestamp 1634918361
transform 1 0 14837 0 1 31343
box 0 0 1 1
use contact_14  contact_14_253
timestamp 1634918361
transform 1 0 14497 0 1 31351
box 0 0 1 1
use contact_13  contact_13_253
timestamp 1634918361
transform 1 0 14501 0 1 31343
box 0 0 1 1
use contact_14  contact_14_254
timestamp 1634918361
transform 1 0 14161 0 1 31351
box 0 0 1 1
use contact_13  contact_13_254
timestamp 1634918361
transform 1 0 14165 0 1 31343
box 0 0 1 1
use contact_7  contact_7_52
timestamp 1634918361
transform 1 0 13821 0 1 31347
box 0 0 1 1
use contact_19  contact_19_190
timestamp 1634918361
transform 1 0 13822 0 1 31352
box 0 0 1 1
use contact_14  contact_14_255
timestamp 1634918361
transform 1 0 13825 0 1 31351
box 0 0 1 1
use contact_13  contact_13_255
timestamp 1634918361
transform 1 0 13829 0 1 31343
box 0 0 1 1
use contact_14  contact_14_256
timestamp 1634918361
transform 1 0 13489 0 1 31351
box 0 0 1 1
use contact_13  contact_13_256
timestamp 1634918361
transform 1 0 13493 0 1 31343
box 0 0 1 1
use contact_14  contact_14_257
timestamp 1634918361
transform 1 0 13153 0 1 31351
box 0 0 1 1
use contact_13  contact_13_257
timestamp 1634918361
transform 1 0 13157 0 1 31343
box 0 0 1 1
use contact_14  contact_14_258
timestamp 1634918361
transform 1 0 12817 0 1 31351
box 0 0 1 1
use contact_13  contact_13_258
timestamp 1634918361
transform 1 0 12821 0 1 31343
box 0 0 1 1
use contact_14  contact_14_259
timestamp 1634918361
transform 1 0 12481 0 1 31351
box 0 0 1 1
use contact_13  contact_13_259
timestamp 1634918361
transform 1 0 12485 0 1 31343
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1634918361
transform 1 0 12141 0 1 31347
box 0 0 1 1
use contact_19  contact_19_191
timestamp 1634918361
transform 1 0 12142 0 1 31352
box 0 0 1 1
use contact_14  contact_14_260
timestamp 1634918361
transform 1 0 12145 0 1 31351
box 0 0 1 1
use contact_13  contact_13_260
timestamp 1634918361
transform 1 0 12149 0 1 31343
box 0 0 1 1
use contact_14  contact_14_261
timestamp 1634918361
transform 1 0 11809 0 1 31351
box 0 0 1 1
use contact_13  contact_13_261
timestamp 1634918361
transform 1 0 11813 0 1 31343
box 0 0 1 1
use contact_14  contact_14_262
timestamp 1634918361
transform 1 0 11473 0 1 31351
box 0 0 1 1
use contact_13  contact_13_262
timestamp 1634918361
transform 1 0 11477 0 1 31343
box 0 0 1 1
use contact_14  contact_14_263
timestamp 1634918361
transform 1 0 11137 0 1 31351
box 0 0 1 1
use contact_13  contact_13_263
timestamp 1634918361
transform 1 0 11141 0 1 31343
box 0 0 1 1
use contact_14  contact_14_264
timestamp 1634918361
transform 1 0 10801 0 1 31351
box 0 0 1 1
use contact_13  contact_13_264
timestamp 1634918361
transform 1 0 10805 0 1 31343
box 0 0 1 1
use contact_7  contact_7_54
timestamp 1634918361
transform 1 0 10461 0 1 31347
box 0 0 1 1
use contact_19  contact_19_192
timestamp 1634918361
transform 1 0 10462 0 1 31352
box 0 0 1 1
use contact_14  contact_14_265
timestamp 1634918361
transform 1 0 10465 0 1 31351
box 0 0 1 1
use contact_13  contact_13_265
timestamp 1634918361
transform 1 0 10469 0 1 31343
box 0 0 1 1
use contact_14  contact_14_266
timestamp 1634918361
transform 1 0 10129 0 1 31351
box 0 0 1 1
use contact_13  contact_13_266
timestamp 1634918361
transform 1 0 10133 0 1 31343
box 0 0 1 1
use contact_14  contact_14_267
timestamp 1634918361
transform 1 0 9793 0 1 31351
box 0 0 1 1
use contact_13  contact_13_267
timestamp 1634918361
transform 1 0 9797 0 1 31343
box 0 0 1 1
use contact_14  contact_14_268
timestamp 1634918361
transform 1 0 9457 0 1 31351
box 0 0 1 1
use contact_13  contact_13_268
timestamp 1634918361
transform 1 0 9461 0 1 31343
box 0 0 1 1
use contact_14  contact_14_269
timestamp 1634918361
transform 1 0 9121 0 1 31351
box 0 0 1 1
use contact_13  contact_13_269
timestamp 1634918361
transform 1 0 9125 0 1 31343
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1634918361
transform 1 0 8781 0 1 31347
box 0 0 1 1
use contact_19  contact_19_193
timestamp 1634918361
transform 1 0 8782 0 1 31352
box 0 0 1 1
use contact_14  contact_14_270
timestamp 1634918361
transform 1 0 8785 0 1 31351
box 0 0 1 1
use contact_13  contact_13_270
timestamp 1634918361
transform 1 0 8789 0 1 31343
box 0 0 1 1
use contact_14  contact_14_271
timestamp 1634918361
transform 1 0 8449 0 1 31351
box 0 0 1 1
use contact_13  contact_13_271
timestamp 1634918361
transform 1 0 8453 0 1 31343
box 0 0 1 1
use contact_14  contact_14_272
timestamp 1634918361
transform 1 0 8113 0 1 31351
box 0 0 1 1
use contact_13  contact_13_272
timestamp 1634918361
transform 1 0 8117 0 1 31343
box 0 0 1 1
use contact_14  contact_14_273
timestamp 1634918361
transform 1 0 7777 0 1 31351
box 0 0 1 1
use contact_13  contact_13_273
timestamp 1634918361
transform 1 0 7781 0 1 31343
box 0 0 1 1
use contact_14  contact_14_274
timestamp 1634918361
transform 1 0 7441 0 1 31351
box 0 0 1 1
use contact_13  contact_13_274
timestamp 1634918361
transform 1 0 7445 0 1 31343
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1634918361
transform 1 0 7101 0 1 31347
box 0 0 1 1
use contact_19  contact_19_194
timestamp 1634918361
transform 1 0 7102 0 1 31352
box 0 0 1 1
use contact_14  contact_14_275
timestamp 1634918361
transform 1 0 7105 0 1 31351
box 0 0 1 1
use contact_13  contact_13_275
timestamp 1634918361
transform 1 0 7109 0 1 31343
box 0 0 1 1
use contact_14  contact_14_276
timestamp 1634918361
transform 1 0 6769 0 1 31351
box 0 0 1 1
use contact_13  contact_13_276
timestamp 1634918361
transform 1 0 6773 0 1 31343
box 0 0 1 1
use contact_14  contact_14_277
timestamp 1634918361
transform 1 0 6433 0 1 31351
box 0 0 1 1
use contact_13  contact_13_277
timestamp 1634918361
transform 1 0 6437 0 1 31343
box 0 0 1 1
use contact_14  contact_14_278
timestamp 1634918361
transform 1 0 6097 0 1 31351
box 0 0 1 1
use contact_13  contact_13_278
timestamp 1634918361
transform 1 0 6101 0 1 31343
box 0 0 1 1
use contact_14  contact_14_279
timestamp 1634918361
transform 1 0 5761 0 1 31351
box 0 0 1 1
use contact_13  contact_13_279
timestamp 1634918361
transform 1 0 5765 0 1 31343
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1634918361
transform 1 0 5421 0 1 31347
box 0 0 1 1
use contact_19  contact_19_195
timestamp 1634918361
transform 1 0 5422 0 1 31352
box 0 0 1 1
use contact_14  contact_14_280
timestamp 1634918361
transform 1 0 5425 0 1 31351
box 0 0 1 1
use contact_13  contact_13_280
timestamp 1634918361
transform 1 0 5429 0 1 31343
box 0 0 1 1
use contact_14  contact_14_281
timestamp 1634918361
transform 1 0 5089 0 1 31351
box 0 0 1 1
use contact_13  contact_13_281
timestamp 1634918361
transform 1 0 5093 0 1 31343
box 0 0 1 1
use contact_14  contact_14_282
timestamp 1634918361
transform 1 0 4753 0 1 31351
box 0 0 1 1
use contact_13  contact_13_282
timestamp 1634918361
transform 1 0 4757 0 1 31343
box 0 0 1 1
use contact_14  contact_14_283
timestamp 1634918361
transform 1 0 4417 0 1 31351
box 0 0 1 1
use contact_13  contact_13_283
timestamp 1634918361
transform 1 0 4421 0 1 31343
box 0 0 1 1
use contact_14  contact_14_284
timestamp 1634918361
transform 1 0 4081 0 1 31351
box 0 0 1 1
use contact_13  contact_13_284
timestamp 1634918361
transform 1 0 4085 0 1 31343
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1634918361
transform 1 0 3741 0 1 31347
box 0 0 1 1
use contact_19  contact_19_196
timestamp 1634918361
transform 1 0 3742 0 1 31352
box 0 0 1 1
use contact_14  contact_14_285
timestamp 1634918361
transform 1 0 3745 0 1 31351
box 0 0 1 1
use contact_13  contact_13_285
timestamp 1634918361
transform 1 0 3749 0 1 31343
box 0 0 1 1
use contact_14  contact_14_286
timestamp 1634918361
transform 1 0 3409 0 1 31351
box 0 0 1 1
use contact_13  contact_13_286
timestamp 1634918361
transform 1 0 3413 0 1 31343
box 0 0 1 1
use contact_14  contact_14_287
timestamp 1634918361
transform 1 0 3073 0 1 31351
box 0 0 1 1
use contact_13  contact_13_287
timestamp 1634918361
transform 1 0 3077 0 1 31343
box 0 0 1 1
use contact_14  contact_14_288
timestamp 1634918361
transform 1 0 2737 0 1 31351
box 0 0 1 1
use contact_13  contact_13_288
timestamp 1634918361
transform 1 0 2741 0 1 31343
box 0 0 1 1
use contact_14  contact_14_289
timestamp 1634918361
transform 1 0 2401 0 1 31351
box 0 0 1 1
use contact_13  contact_13_289
timestamp 1634918361
transform 1 0 2405 0 1 31343
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1634918361
transform 1 0 2061 0 1 31347
box 0 0 1 1
use contact_19  contact_19_197
timestamp 1634918361
transform 1 0 2062 0 1 31352
box 0 0 1 1
use contact_14  contact_14_290
timestamp 1634918361
transform 1 0 2065 0 1 31351
box 0 0 1 1
use contact_13  contact_13_290
timestamp 1634918361
transform 1 0 2069 0 1 31343
box 0 0 1 1
use contact_14  contact_14_291
timestamp 1634918361
transform 1 0 41041 0 1 1727
box 0 0 1 1
use contact_13  contact_13_291
timestamp 1634918361
transform 1 0 41045 0 1 1719
box 0 0 1 1
use contact_7  contact_7_60
timestamp 1634918361
transform 1 0 40701 0 1 1723
box 0 0 1 1
use contact_19  contact_19_198
timestamp 1634918361
transform 1 0 40702 0 1 1728
box 0 0 1 1
use contact_14  contact_14_292
timestamp 1634918361
transform 1 0 40705 0 1 1727
box 0 0 1 1
use contact_13  contact_13_292
timestamp 1634918361
transform 1 0 40709 0 1 1719
box 0 0 1 1
use contact_14  contact_14_293
timestamp 1634918361
transform 1 0 40369 0 1 1727
box 0 0 1 1
use contact_13  contact_13_293
timestamp 1634918361
transform 1 0 40373 0 1 1719
box 0 0 1 1
use contact_14  contact_14_294
timestamp 1634918361
transform 1 0 40033 0 1 1727
box 0 0 1 1
use contact_13  contact_13_294
timestamp 1634918361
transform 1 0 40037 0 1 1719
box 0 0 1 1
use contact_14  contact_14_295
timestamp 1634918361
transform 1 0 39697 0 1 1727
box 0 0 1 1
use contact_13  contact_13_295
timestamp 1634918361
transform 1 0 39701 0 1 1719
box 0 0 1 1
use contact_14  contact_14_296
timestamp 1634918361
transform 1 0 39361 0 1 1727
box 0 0 1 1
use contact_13  contact_13_296
timestamp 1634918361
transform 1 0 39365 0 1 1719
box 0 0 1 1
use contact_7  contact_7_61
timestamp 1634918361
transform 1 0 39021 0 1 1723
box 0 0 1 1
use contact_19  contact_19_199
timestamp 1634918361
transform 1 0 39022 0 1 1728
box 0 0 1 1
use contact_14  contact_14_297
timestamp 1634918361
transform 1 0 39025 0 1 1727
box 0 0 1 1
use contact_13  contact_13_297
timestamp 1634918361
transform 1 0 39029 0 1 1719
box 0 0 1 1
use contact_14  contact_14_298
timestamp 1634918361
transform 1 0 38689 0 1 1727
box 0 0 1 1
use contact_13  contact_13_298
timestamp 1634918361
transform 1 0 38693 0 1 1719
box 0 0 1 1
use contact_14  contact_14_299
timestamp 1634918361
transform 1 0 38353 0 1 1727
box 0 0 1 1
use contact_13  contact_13_299
timestamp 1634918361
transform 1 0 38357 0 1 1719
box 0 0 1 1
use contact_14  contact_14_300
timestamp 1634918361
transform 1 0 38017 0 1 1727
box 0 0 1 1
use contact_13  contact_13_300
timestamp 1634918361
transform 1 0 38021 0 1 1719
box 0 0 1 1
use contact_14  contact_14_301
timestamp 1634918361
transform 1 0 37681 0 1 1727
box 0 0 1 1
use contact_13  contact_13_301
timestamp 1634918361
transform 1 0 37685 0 1 1719
box 0 0 1 1
use contact_7  contact_7_62
timestamp 1634918361
transform 1 0 37341 0 1 1723
box 0 0 1 1
use contact_19  contact_19_200
timestamp 1634918361
transform 1 0 37342 0 1 1728
box 0 0 1 1
use contact_14  contact_14_302
timestamp 1634918361
transform 1 0 37345 0 1 1727
box 0 0 1 1
use contact_13  contact_13_302
timestamp 1634918361
transform 1 0 37349 0 1 1719
box 0 0 1 1
use contact_14  contact_14_303
timestamp 1634918361
transform 1 0 37009 0 1 1727
box 0 0 1 1
use contact_13  contact_13_303
timestamp 1634918361
transform 1 0 37013 0 1 1719
box 0 0 1 1
use contact_14  contact_14_304
timestamp 1634918361
transform 1 0 36673 0 1 1727
box 0 0 1 1
use contact_13  contact_13_304
timestamp 1634918361
transform 1 0 36677 0 1 1719
box 0 0 1 1
use contact_14  contact_14_305
timestamp 1634918361
transform 1 0 36337 0 1 1727
box 0 0 1 1
use contact_13  contact_13_305
timestamp 1634918361
transform 1 0 36341 0 1 1719
box 0 0 1 1
use contact_14  contact_14_306
timestamp 1634918361
transform 1 0 36001 0 1 1727
box 0 0 1 1
use contact_13  contact_13_306
timestamp 1634918361
transform 1 0 36005 0 1 1719
box 0 0 1 1
use contact_7  contact_7_63
timestamp 1634918361
transform 1 0 35661 0 1 1723
box 0 0 1 1
use contact_19  contact_19_201
timestamp 1634918361
transform 1 0 35662 0 1 1728
box 0 0 1 1
use contact_14  contact_14_307
timestamp 1634918361
transform 1 0 35665 0 1 1727
box 0 0 1 1
use contact_13  contact_13_307
timestamp 1634918361
transform 1 0 35669 0 1 1719
box 0 0 1 1
use contact_14  contact_14_308
timestamp 1634918361
transform 1 0 35329 0 1 1727
box 0 0 1 1
use contact_13  contact_13_308
timestamp 1634918361
transform 1 0 35333 0 1 1719
box 0 0 1 1
use contact_14  contact_14_309
timestamp 1634918361
transform 1 0 34993 0 1 1727
box 0 0 1 1
use contact_13  contact_13_309
timestamp 1634918361
transform 1 0 34997 0 1 1719
box 0 0 1 1
use contact_14  contact_14_310
timestamp 1634918361
transform 1 0 34657 0 1 1727
box 0 0 1 1
use contact_13  contact_13_310
timestamp 1634918361
transform 1 0 34661 0 1 1719
box 0 0 1 1
use contact_14  contact_14_311
timestamp 1634918361
transform 1 0 34321 0 1 1727
box 0 0 1 1
use contact_13  contact_13_311
timestamp 1634918361
transform 1 0 34325 0 1 1719
box 0 0 1 1
use contact_7  contact_7_64
timestamp 1634918361
transform 1 0 33981 0 1 1723
box 0 0 1 1
use contact_19  contact_19_202
timestamp 1634918361
transform 1 0 33982 0 1 1728
box 0 0 1 1
use contact_14  contact_14_312
timestamp 1634918361
transform 1 0 33985 0 1 1727
box 0 0 1 1
use contact_13  contact_13_312
timestamp 1634918361
transform 1 0 33989 0 1 1719
box 0 0 1 1
use contact_14  contact_14_313
timestamp 1634918361
transform 1 0 33649 0 1 1727
box 0 0 1 1
use contact_13  contact_13_313
timestamp 1634918361
transform 1 0 33653 0 1 1719
box 0 0 1 1
use contact_14  contact_14_314
timestamp 1634918361
transform 1 0 33313 0 1 1727
box 0 0 1 1
use contact_13  contact_13_314
timestamp 1634918361
transform 1 0 33317 0 1 1719
box 0 0 1 1
use contact_14  contact_14_315
timestamp 1634918361
transform 1 0 32977 0 1 1727
box 0 0 1 1
use contact_13  contact_13_315
timestamp 1634918361
transform 1 0 32981 0 1 1719
box 0 0 1 1
use contact_14  contact_14_316
timestamp 1634918361
transform 1 0 32641 0 1 1727
box 0 0 1 1
use contact_13  contact_13_316
timestamp 1634918361
transform 1 0 32645 0 1 1719
box 0 0 1 1
use contact_7  contact_7_65
timestamp 1634918361
transform 1 0 32301 0 1 1723
box 0 0 1 1
use contact_19  contact_19_203
timestamp 1634918361
transform 1 0 32302 0 1 1728
box 0 0 1 1
use contact_14  contact_14_317
timestamp 1634918361
transform 1 0 32305 0 1 1727
box 0 0 1 1
use contact_13  contact_13_317
timestamp 1634918361
transform 1 0 32309 0 1 1719
box 0 0 1 1
use contact_14  contact_14_318
timestamp 1634918361
transform 1 0 31969 0 1 1727
box 0 0 1 1
use contact_13  contact_13_318
timestamp 1634918361
transform 1 0 31973 0 1 1719
box 0 0 1 1
use contact_14  contact_14_319
timestamp 1634918361
transform 1 0 31633 0 1 1727
box 0 0 1 1
use contact_13  contact_13_319
timestamp 1634918361
transform 1 0 31637 0 1 1719
box 0 0 1 1
use contact_14  contact_14_320
timestamp 1634918361
transform 1 0 31297 0 1 1727
box 0 0 1 1
use contact_13  contact_13_320
timestamp 1634918361
transform 1 0 31301 0 1 1719
box 0 0 1 1
use contact_14  contact_14_321
timestamp 1634918361
transform 1 0 30961 0 1 1727
box 0 0 1 1
use contact_13  contact_13_321
timestamp 1634918361
transform 1 0 30965 0 1 1719
box 0 0 1 1
use contact_7  contact_7_66
timestamp 1634918361
transform 1 0 30621 0 1 1723
box 0 0 1 1
use contact_19  contact_19_204
timestamp 1634918361
transform 1 0 30622 0 1 1728
box 0 0 1 1
use contact_14  contact_14_322
timestamp 1634918361
transform 1 0 30625 0 1 1727
box 0 0 1 1
use contact_13  contact_13_322
timestamp 1634918361
transform 1 0 30629 0 1 1719
box 0 0 1 1
use contact_14  contact_14_323
timestamp 1634918361
transform 1 0 30289 0 1 1727
box 0 0 1 1
use contact_13  contact_13_323
timestamp 1634918361
transform 1 0 30293 0 1 1719
box 0 0 1 1
use contact_14  contact_14_324
timestamp 1634918361
transform 1 0 29953 0 1 1727
box 0 0 1 1
use contact_13  contact_13_324
timestamp 1634918361
transform 1 0 29957 0 1 1719
box 0 0 1 1
use contact_14  contact_14_325
timestamp 1634918361
transform 1 0 29617 0 1 1727
box 0 0 1 1
use contact_13  contact_13_325
timestamp 1634918361
transform 1 0 29621 0 1 1719
box 0 0 1 1
use contact_14  contact_14_326
timestamp 1634918361
transform 1 0 29281 0 1 1727
box 0 0 1 1
use contact_13  contact_13_326
timestamp 1634918361
transform 1 0 29285 0 1 1719
box 0 0 1 1
use contact_7  contact_7_67
timestamp 1634918361
transform 1 0 28941 0 1 1723
box 0 0 1 1
use contact_19  contact_19_205
timestamp 1634918361
transform 1 0 28942 0 1 1728
box 0 0 1 1
use contact_14  contact_14_327
timestamp 1634918361
transform 1 0 28945 0 1 1727
box 0 0 1 1
use contact_13  contact_13_327
timestamp 1634918361
transform 1 0 28949 0 1 1719
box 0 0 1 1
use contact_14  contact_14_328
timestamp 1634918361
transform 1 0 28609 0 1 1727
box 0 0 1 1
use contact_13  contact_13_328
timestamp 1634918361
transform 1 0 28613 0 1 1719
box 0 0 1 1
use contact_14  contact_14_329
timestamp 1634918361
transform 1 0 28273 0 1 1727
box 0 0 1 1
use contact_13  contact_13_329
timestamp 1634918361
transform 1 0 28277 0 1 1719
box 0 0 1 1
use contact_14  contact_14_330
timestamp 1634918361
transform 1 0 27937 0 1 1727
box 0 0 1 1
use contact_13  contact_13_330
timestamp 1634918361
transform 1 0 27941 0 1 1719
box 0 0 1 1
use contact_14  contact_14_331
timestamp 1634918361
transform 1 0 27601 0 1 1727
box 0 0 1 1
use contact_13  contact_13_331
timestamp 1634918361
transform 1 0 27605 0 1 1719
box 0 0 1 1
use contact_7  contact_7_68
timestamp 1634918361
transform 1 0 27261 0 1 1723
box 0 0 1 1
use contact_19  contact_19_206
timestamp 1634918361
transform 1 0 27262 0 1 1728
box 0 0 1 1
use contact_14  contact_14_332
timestamp 1634918361
transform 1 0 27265 0 1 1727
box 0 0 1 1
use contact_13  contact_13_332
timestamp 1634918361
transform 1 0 27269 0 1 1719
box 0 0 1 1
use contact_14  contact_14_333
timestamp 1634918361
transform 1 0 26929 0 1 1727
box 0 0 1 1
use contact_13  contact_13_333
timestamp 1634918361
transform 1 0 26933 0 1 1719
box 0 0 1 1
use contact_14  contact_14_334
timestamp 1634918361
transform 1 0 26593 0 1 1727
box 0 0 1 1
use contact_13  contact_13_334
timestamp 1634918361
transform 1 0 26597 0 1 1719
box 0 0 1 1
use contact_14  contact_14_335
timestamp 1634918361
transform 1 0 26257 0 1 1727
box 0 0 1 1
use contact_13  contact_13_335
timestamp 1634918361
transform 1 0 26261 0 1 1719
box 0 0 1 1
use contact_14  contact_14_336
timestamp 1634918361
transform 1 0 25921 0 1 1727
box 0 0 1 1
use contact_13  contact_13_336
timestamp 1634918361
transform 1 0 25925 0 1 1719
box 0 0 1 1
use contact_7  contact_7_69
timestamp 1634918361
transform 1 0 25581 0 1 1723
box 0 0 1 1
use contact_19  contact_19_207
timestamp 1634918361
transform 1 0 25582 0 1 1728
box 0 0 1 1
use contact_14  contact_14_337
timestamp 1634918361
transform 1 0 25585 0 1 1727
box 0 0 1 1
use contact_13  contact_13_337
timestamp 1634918361
transform 1 0 25589 0 1 1719
box 0 0 1 1
use contact_14  contact_14_338
timestamp 1634918361
transform 1 0 25249 0 1 1727
box 0 0 1 1
use contact_13  contact_13_338
timestamp 1634918361
transform 1 0 25253 0 1 1719
box 0 0 1 1
use contact_14  contact_14_339
timestamp 1634918361
transform 1 0 24913 0 1 1727
box 0 0 1 1
use contact_13  contact_13_339
timestamp 1634918361
transform 1 0 24917 0 1 1719
box 0 0 1 1
use contact_14  contact_14_340
timestamp 1634918361
transform 1 0 24577 0 1 1727
box 0 0 1 1
use contact_13  contact_13_340
timestamp 1634918361
transform 1 0 24581 0 1 1719
box 0 0 1 1
use contact_14  contact_14_341
timestamp 1634918361
transform 1 0 24241 0 1 1727
box 0 0 1 1
use contact_13  contact_13_341
timestamp 1634918361
transform 1 0 24245 0 1 1719
box 0 0 1 1
use contact_7  contact_7_70
timestamp 1634918361
transform 1 0 23901 0 1 1723
box 0 0 1 1
use contact_19  contact_19_208
timestamp 1634918361
transform 1 0 23902 0 1 1728
box 0 0 1 1
use contact_14  contact_14_342
timestamp 1634918361
transform 1 0 23905 0 1 1727
box 0 0 1 1
use contact_13  contact_13_342
timestamp 1634918361
transform 1 0 23909 0 1 1719
box 0 0 1 1
use contact_14  contact_14_343
timestamp 1634918361
transform 1 0 23569 0 1 1727
box 0 0 1 1
use contact_13  contact_13_343
timestamp 1634918361
transform 1 0 23573 0 1 1719
box 0 0 1 1
use contact_14  contact_14_344
timestamp 1634918361
transform 1 0 23233 0 1 1727
box 0 0 1 1
use contact_13  contact_13_344
timestamp 1634918361
transform 1 0 23237 0 1 1719
box 0 0 1 1
use contact_14  contact_14_345
timestamp 1634918361
transform 1 0 22897 0 1 1727
box 0 0 1 1
use contact_13  contact_13_345
timestamp 1634918361
transform 1 0 22901 0 1 1719
box 0 0 1 1
use contact_14  contact_14_346
timestamp 1634918361
transform 1 0 22561 0 1 1727
box 0 0 1 1
use contact_13  contact_13_346
timestamp 1634918361
transform 1 0 22565 0 1 1719
box 0 0 1 1
use contact_7  contact_7_71
timestamp 1634918361
transform 1 0 22221 0 1 1723
box 0 0 1 1
use contact_19  contact_19_209
timestamp 1634918361
transform 1 0 22222 0 1 1728
box 0 0 1 1
use contact_14  contact_14_347
timestamp 1634918361
transform 1 0 22225 0 1 1727
box 0 0 1 1
use contact_13  contact_13_347
timestamp 1634918361
transform 1 0 22229 0 1 1719
box 0 0 1 1
use contact_14  contact_14_348
timestamp 1634918361
transform 1 0 21889 0 1 1727
box 0 0 1 1
use contact_13  contact_13_348
timestamp 1634918361
transform 1 0 21893 0 1 1719
box 0 0 1 1
use contact_14  contact_14_349
timestamp 1634918361
transform 1 0 21553 0 1 1727
box 0 0 1 1
use contact_13  contact_13_349
timestamp 1634918361
transform 1 0 21557 0 1 1719
box 0 0 1 1
use contact_14  contact_14_350
timestamp 1634918361
transform 1 0 21217 0 1 1727
box 0 0 1 1
use contact_13  contact_13_350
timestamp 1634918361
transform 1 0 21221 0 1 1719
box 0 0 1 1
use contact_14  contact_14_351
timestamp 1634918361
transform 1 0 20881 0 1 1727
box 0 0 1 1
use contact_13  contact_13_351
timestamp 1634918361
transform 1 0 20885 0 1 1719
box 0 0 1 1
use contact_7  contact_7_72
timestamp 1634918361
transform 1 0 20541 0 1 1723
box 0 0 1 1
use contact_19  contact_19_210
timestamp 1634918361
transform 1 0 20542 0 1 1728
box 0 0 1 1
use contact_14  contact_14_352
timestamp 1634918361
transform 1 0 20545 0 1 1727
box 0 0 1 1
use contact_13  contact_13_352
timestamp 1634918361
transform 1 0 20549 0 1 1719
box 0 0 1 1
use contact_14  contact_14_353
timestamp 1634918361
transform 1 0 20209 0 1 1727
box 0 0 1 1
use contact_13  contact_13_353
timestamp 1634918361
transform 1 0 20213 0 1 1719
box 0 0 1 1
use contact_14  contact_14_354
timestamp 1634918361
transform 1 0 19873 0 1 1727
box 0 0 1 1
use contact_13  contact_13_354
timestamp 1634918361
transform 1 0 19877 0 1 1719
box 0 0 1 1
use contact_14  contact_14_355
timestamp 1634918361
transform 1 0 19537 0 1 1727
box 0 0 1 1
use contact_13  contact_13_355
timestamp 1634918361
transform 1 0 19541 0 1 1719
box 0 0 1 1
use contact_14  contact_14_356
timestamp 1634918361
transform 1 0 19201 0 1 1727
box 0 0 1 1
use contact_13  contact_13_356
timestamp 1634918361
transform 1 0 19205 0 1 1719
box 0 0 1 1
use contact_7  contact_7_73
timestamp 1634918361
transform 1 0 18861 0 1 1723
box 0 0 1 1
use contact_19  contact_19_211
timestamp 1634918361
transform 1 0 18862 0 1 1728
box 0 0 1 1
use contact_14  contact_14_357
timestamp 1634918361
transform 1 0 18865 0 1 1727
box 0 0 1 1
use contact_13  contact_13_357
timestamp 1634918361
transform 1 0 18869 0 1 1719
box 0 0 1 1
use contact_14  contact_14_358
timestamp 1634918361
transform 1 0 18529 0 1 1727
box 0 0 1 1
use contact_13  contact_13_358
timestamp 1634918361
transform 1 0 18533 0 1 1719
box 0 0 1 1
use contact_14  contact_14_359
timestamp 1634918361
transform 1 0 18193 0 1 1727
box 0 0 1 1
use contact_13  contact_13_359
timestamp 1634918361
transform 1 0 18197 0 1 1719
box 0 0 1 1
use contact_14  contact_14_360
timestamp 1634918361
transform 1 0 17857 0 1 1727
box 0 0 1 1
use contact_13  contact_13_360
timestamp 1634918361
transform 1 0 17861 0 1 1719
box 0 0 1 1
use contact_14  contact_14_361
timestamp 1634918361
transform 1 0 17521 0 1 1727
box 0 0 1 1
use contact_13  contact_13_361
timestamp 1634918361
transform 1 0 17525 0 1 1719
box 0 0 1 1
use contact_7  contact_7_74
timestamp 1634918361
transform 1 0 17181 0 1 1723
box 0 0 1 1
use contact_19  contact_19_212
timestamp 1634918361
transform 1 0 17182 0 1 1728
box 0 0 1 1
use contact_14  contact_14_362
timestamp 1634918361
transform 1 0 17185 0 1 1727
box 0 0 1 1
use contact_13  contact_13_362
timestamp 1634918361
transform 1 0 17189 0 1 1719
box 0 0 1 1
use contact_14  contact_14_363
timestamp 1634918361
transform 1 0 16849 0 1 1727
box 0 0 1 1
use contact_13  contact_13_363
timestamp 1634918361
transform 1 0 16853 0 1 1719
box 0 0 1 1
use contact_14  contact_14_364
timestamp 1634918361
transform 1 0 16513 0 1 1727
box 0 0 1 1
use contact_13  contact_13_364
timestamp 1634918361
transform 1 0 16517 0 1 1719
box 0 0 1 1
use contact_14  contact_14_365
timestamp 1634918361
transform 1 0 16177 0 1 1727
box 0 0 1 1
use contact_13  contact_13_365
timestamp 1634918361
transform 1 0 16181 0 1 1719
box 0 0 1 1
use contact_14  contact_14_366
timestamp 1634918361
transform 1 0 15841 0 1 1727
box 0 0 1 1
use contact_13  contact_13_366
timestamp 1634918361
transform 1 0 15845 0 1 1719
box 0 0 1 1
use contact_7  contact_7_75
timestamp 1634918361
transform 1 0 15501 0 1 1723
box 0 0 1 1
use contact_19  contact_19_213
timestamp 1634918361
transform 1 0 15502 0 1 1728
box 0 0 1 1
use contact_14  contact_14_367
timestamp 1634918361
transform 1 0 15505 0 1 1727
box 0 0 1 1
use contact_13  contact_13_367
timestamp 1634918361
transform 1 0 15509 0 1 1719
box 0 0 1 1
use contact_14  contact_14_368
timestamp 1634918361
transform 1 0 15169 0 1 1727
box 0 0 1 1
use contact_13  contact_13_368
timestamp 1634918361
transform 1 0 15173 0 1 1719
box 0 0 1 1
use contact_14  contact_14_369
timestamp 1634918361
transform 1 0 14833 0 1 1727
box 0 0 1 1
use contact_13  contact_13_369
timestamp 1634918361
transform 1 0 14837 0 1 1719
box 0 0 1 1
use contact_14  contact_14_370
timestamp 1634918361
transform 1 0 14497 0 1 1727
box 0 0 1 1
use contact_13  contact_13_370
timestamp 1634918361
transform 1 0 14501 0 1 1719
box 0 0 1 1
use contact_14  contact_14_371
timestamp 1634918361
transform 1 0 14161 0 1 1727
box 0 0 1 1
use contact_13  contact_13_371
timestamp 1634918361
transform 1 0 14165 0 1 1719
box 0 0 1 1
use contact_7  contact_7_76
timestamp 1634918361
transform 1 0 13821 0 1 1723
box 0 0 1 1
use contact_19  contact_19_214
timestamp 1634918361
transform 1 0 13822 0 1 1728
box 0 0 1 1
use contact_14  contact_14_372
timestamp 1634918361
transform 1 0 13825 0 1 1727
box 0 0 1 1
use contact_13  contact_13_372
timestamp 1634918361
transform 1 0 13829 0 1 1719
box 0 0 1 1
use contact_14  contact_14_373
timestamp 1634918361
transform 1 0 13489 0 1 1727
box 0 0 1 1
use contact_13  contact_13_373
timestamp 1634918361
transform 1 0 13493 0 1 1719
box 0 0 1 1
use contact_14  contact_14_374
timestamp 1634918361
transform 1 0 13153 0 1 1727
box 0 0 1 1
use contact_13  contact_13_374
timestamp 1634918361
transform 1 0 13157 0 1 1719
box 0 0 1 1
use contact_14  contact_14_375
timestamp 1634918361
transform 1 0 12817 0 1 1727
box 0 0 1 1
use contact_13  contact_13_375
timestamp 1634918361
transform 1 0 12821 0 1 1719
box 0 0 1 1
use contact_14  contact_14_376
timestamp 1634918361
transform 1 0 12481 0 1 1727
box 0 0 1 1
use contact_13  contact_13_376
timestamp 1634918361
transform 1 0 12485 0 1 1719
box 0 0 1 1
use contact_7  contact_7_77
timestamp 1634918361
transform 1 0 12141 0 1 1723
box 0 0 1 1
use contact_19  contact_19_215
timestamp 1634918361
transform 1 0 12142 0 1 1728
box 0 0 1 1
use contact_14  contact_14_377
timestamp 1634918361
transform 1 0 12145 0 1 1727
box 0 0 1 1
use contact_13  contact_13_377
timestamp 1634918361
transform 1 0 12149 0 1 1719
box 0 0 1 1
use contact_14  contact_14_378
timestamp 1634918361
transform 1 0 11809 0 1 1727
box 0 0 1 1
use contact_13  contact_13_378
timestamp 1634918361
transform 1 0 11813 0 1 1719
box 0 0 1 1
use contact_14  contact_14_379
timestamp 1634918361
transform 1 0 11473 0 1 1727
box 0 0 1 1
use contact_13  contact_13_379
timestamp 1634918361
transform 1 0 11477 0 1 1719
box 0 0 1 1
use contact_14  contact_14_380
timestamp 1634918361
transform 1 0 11137 0 1 1727
box 0 0 1 1
use contact_13  contact_13_380
timestamp 1634918361
transform 1 0 11141 0 1 1719
box 0 0 1 1
use contact_14  contact_14_381
timestamp 1634918361
transform 1 0 10801 0 1 1727
box 0 0 1 1
use contact_13  contact_13_381
timestamp 1634918361
transform 1 0 10805 0 1 1719
box 0 0 1 1
use contact_7  contact_7_78
timestamp 1634918361
transform 1 0 10461 0 1 1723
box 0 0 1 1
use contact_19  contact_19_216
timestamp 1634918361
transform 1 0 10462 0 1 1728
box 0 0 1 1
use contact_14  contact_14_382
timestamp 1634918361
transform 1 0 10465 0 1 1727
box 0 0 1 1
use contact_13  contact_13_382
timestamp 1634918361
transform 1 0 10469 0 1 1719
box 0 0 1 1
use contact_14  contact_14_383
timestamp 1634918361
transform 1 0 10129 0 1 1727
box 0 0 1 1
use contact_13  contact_13_383
timestamp 1634918361
transform 1 0 10133 0 1 1719
box 0 0 1 1
use contact_14  contact_14_384
timestamp 1634918361
transform 1 0 9793 0 1 1727
box 0 0 1 1
use contact_13  contact_13_384
timestamp 1634918361
transform 1 0 9797 0 1 1719
box 0 0 1 1
use contact_14  contact_14_385
timestamp 1634918361
transform 1 0 9457 0 1 1727
box 0 0 1 1
use contact_13  contact_13_385
timestamp 1634918361
transform 1 0 9461 0 1 1719
box 0 0 1 1
use contact_14  contact_14_386
timestamp 1634918361
transform 1 0 9121 0 1 1727
box 0 0 1 1
use contact_13  contact_13_386
timestamp 1634918361
transform 1 0 9125 0 1 1719
box 0 0 1 1
use contact_7  contact_7_79
timestamp 1634918361
transform 1 0 8781 0 1 1723
box 0 0 1 1
use contact_19  contact_19_217
timestamp 1634918361
transform 1 0 8782 0 1 1728
box 0 0 1 1
use contact_14  contact_14_387
timestamp 1634918361
transform 1 0 8785 0 1 1727
box 0 0 1 1
use contact_13  contact_13_387
timestamp 1634918361
transform 1 0 8789 0 1 1719
box 0 0 1 1
use contact_14  contact_14_388
timestamp 1634918361
transform 1 0 8449 0 1 1727
box 0 0 1 1
use contact_13  contact_13_388
timestamp 1634918361
transform 1 0 8453 0 1 1719
box 0 0 1 1
use contact_14  contact_14_389
timestamp 1634918361
transform 1 0 8113 0 1 1727
box 0 0 1 1
use contact_13  contact_13_389
timestamp 1634918361
transform 1 0 8117 0 1 1719
box 0 0 1 1
use contact_14  contact_14_390
timestamp 1634918361
transform 1 0 7777 0 1 1727
box 0 0 1 1
use contact_13  contact_13_390
timestamp 1634918361
transform 1 0 7781 0 1 1719
box 0 0 1 1
use contact_14  contact_14_391
timestamp 1634918361
transform 1 0 7441 0 1 1727
box 0 0 1 1
use contact_13  contact_13_391
timestamp 1634918361
transform 1 0 7445 0 1 1719
box 0 0 1 1
use contact_7  contact_7_80
timestamp 1634918361
transform 1 0 7101 0 1 1723
box 0 0 1 1
use contact_19  contact_19_218
timestamp 1634918361
transform 1 0 7102 0 1 1728
box 0 0 1 1
use contact_14  contact_14_392
timestamp 1634918361
transform 1 0 7105 0 1 1727
box 0 0 1 1
use contact_13  contact_13_392
timestamp 1634918361
transform 1 0 7109 0 1 1719
box 0 0 1 1
use contact_14  contact_14_393
timestamp 1634918361
transform 1 0 6769 0 1 1727
box 0 0 1 1
use contact_13  contact_13_393
timestamp 1634918361
transform 1 0 6773 0 1 1719
box 0 0 1 1
use contact_14  contact_14_394
timestamp 1634918361
transform 1 0 6433 0 1 1727
box 0 0 1 1
use contact_13  contact_13_394
timestamp 1634918361
transform 1 0 6437 0 1 1719
box 0 0 1 1
use contact_14  contact_14_395
timestamp 1634918361
transform 1 0 6097 0 1 1727
box 0 0 1 1
use contact_13  contact_13_395
timestamp 1634918361
transform 1 0 6101 0 1 1719
box 0 0 1 1
use contact_14  contact_14_396
timestamp 1634918361
transform 1 0 5761 0 1 1727
box 0 0 1 1
use contact_13  contact_13_396
timestamp 1634918361
transform 1 0 5765 0 1 1719
box 0 0 1 1
use contact_7  contact_7_81
timestamp 1634918361
transform 1 0 5421 0 1 1723
box 0 0 1 1
use contact_19  contact_19_219
timestamp 1634918361
transform 1 0 5422 0 1 1728
box 0 0 1 1
use contact_14  contact_14_397
timestamp 1634918361
transform 1 0 5425 0 1 1727
box 0 0 1 1
use contact_13  contact_13_397
timestamp 1634918361
transform 1 0 5429 0 1 1719
box 0 0 1 1
use contact_14  contact_14_398
timestamp 1634918361
transform 1 0 5089 0 1 1727
box 0 0 1 1
use contact_13  contact_13_398
timestamp 1634918361
transform 1 0 5093 0 1 1719
box 0 0 1 1
use contact_14  contact_14_399
timestamp 1634918361
transform 1 0 4753 0 1 1727
box 0 0 1 1
use contact_13  contact_13_399
timestamp 1634918361
transform 1 0 4757 0 1 1719
box 0 0 1 1
use contact_14  contact_14_400
timestamp 1634918361
transform 1 0 4417 0 1 1727
box 0 0 1 1
use contact_13  contact_13_400
timestamp 1634918361
transform 1 0 4421 0 1 1719
box 0 0 1 1
use contact_14  contact_14_401
timestamp 1634918361
transform 1 0 4081 0 1 1727
box 0 0 1 1
use contact_13  contact_13_401
timestamp 1634918361
transform 1 0 4085 0 1 1719
box 0 0 1 1
use contact_7  contact_7_82
timestamp 1634918361
transform 1 0 3741 0 1 1723
box 0 0 1 1
use contact_19  contact_19_220
timestamp 1634918361
transform 1 0 3742 0 1 1728
box 0 0 1 1
use contact_14  contact_14_402
timestamp 1634918361
transform 1 0 3745 0 1 1727
box 0 0 1 1
use contact_13  contact_13_402
timestamp 1634918361
transform 1 0 3749 0 1 1719
box 0 0 1 1
use contact_14  contact_14_403
timestamp 1634918361
transform 1 0 3409 0 1 1727
box 0 0 1 1
use contact_13  contact_13_403
timestamp 1634918361
transform 1 0 3413 0 1 1719
box 0 0 1 1
use contact_14  contact_14_404
timestamp 1634918361
transform 1 0 3073 0 1 1727
box 0 0 1 1
use contact_13  contact_13_404
timestamp 1634918361
transform 1 0 3077 0 1 1719
box 0 0 1 1
use contact_14  contact_14_405
timestamp 1634918361
transform 1 0 2737 0 1 1727
box 0 0 1 1
use contact_13  contact_13_405
timestamp 1634918361
transform 1 0 2741 0 1 1719
box 0 0 1 1
use contact_14  contact_14_406
timestamp 1634918361
transform 1 0 2401 0 1 1727
box 0 0 1 1
use contact_13  contact_13_406
timestamp 1634918361
transform 1 0 2405 0 1 1719
box 0 0 1 1
use contact_7  contact_7_83
timestamp 1634918361
transform 1 0 2061 0 1 1723
box 0 0 1 1
use contact_19  contact_19_221
timestamp 1634918361
transform 1 0 2062 0 1 1728
box 0 0 1 1
use contact_14  contact_14_407
timestamp 1634918361
transform 1 0 2065 0 1 1727
box 0 0 1 1
use contact_13  contact_13_407
timestamp 1634918361
transform 1 0 2069 0 1 1719
box 0 0 1 1
use contact_7  contact_7_84
timestamp 1634918361
transform 1 0 35129 0 1 9697
box 0 0 1 1
use contact_7  contact_7_85
timestamp 1634918361
transform 1 0 35129 0 1 11397
box 0 0 1 1
use contact_7  contact_7_86
timestamp 1634918361
transform 1 0 35129 0 1 12525
box 0 0 1 1
use contact_7  contact_7_87
timestamp 1634918361
transform 1 0 35129 0 1 14225
box 0 0 1 1
use contact_7  contact_7_88
timestamp 1634918361
transform 1 0 24139 0 1 25286
box 0 0 1 1
use contact_19  contact_19_222
timestamp 1634918361
transform 1 0 24140 0 1 25291
box 0 0 1 1
use contact_7  contact_7_89
timestamp 1634918361
transform 1 0 23145 0 1 25286
box 0 0 1 1
use contact_19  contact_19_223
timestamp 1634918361
transform 1 0 23146 0 1 25291
box 0 0 1 1
use contact_7  contact_7_90
timestamp 1634918361
transform 1 0 22891 0 1 25286
box 0 0 1 1
use contact_19  contact_19_224
timestamp 1634918361
transform 1 0 22892 0 1 25291
box 0 0 1 1
use contact_7  contact_7_91
timestamp 1634918361
transform 1 0 21897 0 1 25286
box 0 0 1 1
use contact_19  contact_19_225
timestamp 1634918361
transform 1 0 21898 0 1 25291
box 0 0 1 1
use contact_7  contact_7_92
timestamp 1634918361
transform 1 0 21643 0 1 25286
box 0 0 1 1
use contact_19  contact_19_226
timestamp 1634918361
transform 1 0 21644 0 1 25291
box 0 0 1 1
use contact_7  contact_7_93
timestamp 1634918361
transform 1 0 20649 0 1 25286
box 0 0 1 1
use contact_19  contact_19_227
timestamp 1634918361
transform 1 0 20650 0 1 25291
box 0 0 1 1
use contact_7  contact_7_94
timestamp 1634918361
transform 1 0 20395 0 1 25286
box 0 0 1 1
use contact_19  contact_19_228
timestamp 1634918361
transform 1 0 20396 0 1 25291
box 0 0 1 1
use contact_7  contact_7_95
timestamp 1634918361
transform 1 0 19401 0 1 25286
box 0 0 1 1
use contact_19  contact_19_229
timestamp 1634918361
transform 1 0 19402 0 1 25291
box 0 0 1 1
use contact_7  contact_7_96
timestamp 1634918361
transform 1 0 37442 0 1 29838
box 0 0 1 1
use contact_7  contact_7_97
timestamp 1634918361
transform 1 0 40579 0 1 29943
box 0 0 1 1
use contact_7  contact_7_98
timestamp 1634918361
transform 1 0 14335 0 1 3127
box 0 0 1 1
use contact_7  contact_7_99
timestamp 1634918361
transform 1 0 13167 0 1 3127
box 0 0 1 1
use contact_7  contact_7_100
timestamp 1634918361
transform 1 0 11999 0 1 3127
box 0 0 1 1
use contact_7  contact_7_101
timestamp 1634918361
transform 1 0 10831 0 1 3127
box 0 0 1 1
use contact_7  contact_7_102
timestamp 1634918361
transform 1 0 8495 0 1 26197
box 0 0 1 1
use contact_7  contact_7_103
timestamp 1634918361
transform 1 0 8495 0 1 24497
box 0 0 1 1
use contact_7  contact_7_104
timestamp 1634918361
transform 1 0 8495 0 1 23369
box 0 0 1 1
use contact_7  contact_7_105
timestamp 1634918361
transform 1 0 8495 0 1 21669
box 0 0 1 1
use contact_7  contact_7_106
timestamp 1634918361
transform 1 0 24139 0 1 10612
box 0 0 1 1
use contact_19  contact_19_230
timestamp 1634918361
transform 1 0 24140 0 1 10617
box 0 0 1 1
use contact_7  contact_7_107
timestamp 1634918361
transform 1 0 23145 0 1 10612
box 0 0 1 1
use contact_19  contact_19_231
timestamp 1634918361
transform 1 0 23146 0 1 10617
box 0 0 1 1
use contact_7  contact_7_108
timestamp 1634918361
transform 1 0 22891 0 1 10612
box 0 0 1 1
use contact_19  contact_19_232
timestamp 1634918361
transform 1 0 22892 0 1 10617
box 0 0 1 1
use contact_7  contact_7_109
timestamp 1634918361
transform 1 0 21897 0 1 10612
box 0 0 1 1
use contact_19  contact_19_233
timestamp 1634918361
transform 1 0 21898 0 1 10617
box 0 0 1 1
use contact_7  contact_7_110
timestamp 1634918361
transform 1 0 21643 0 1 10612
box 0 0 1 1
use contact_19  contact_19_234
timestamp 1634918361
transform 1 0 21644 0 1 10617
box 0 0 1 1
use contact_7  contact_7_111
timestamp 1634918361
transform 1 0 20649 0 1 10612
box 0 0 1 1
use contact_19  contact_19_235
timestamp 1634918361
transform 1 0 20650 0 1 10617
box 0 0 1 1
use contact_7  contact_7_112
timestamp 1634918361
transform 1 0 20395 0 1 10612
box 0 0 1 1
use contact_19  contact_19_236
timestamp 1634918361
transform 1 0 20396 0 1 10617
box 0 0 1 1
use contact_7  contact_7_113
timestamp 1634918361
transform 1 0 19401 0 1 10612
box 0 0 1 1
use contact_19  contact_19_237
timestamp 1634918361
transform 1 0 19402 0 1 10617
box 0 0 1 1
use contact_7  contact_7_114
timestamp 1634918361
transform 1 0 23679 0 1 3127
box 0 0 1 1
use contact_7  contact_7_115
timestamp 1634918361
transform 1 0 22511 0 1 3127
box 0 0 1 1
use contact_7  contact_7_116
timestamp 1634918361
transform 1 0 21343 0 1 3127
box 0 0 1 1
use contact_7  contact_7_117
timestamp 1634918361
transform 1 0 20175 0 1 3127
box 0 0 1 1
use contact_7  contact_7_118
timestamp 1634918361
transform 1 0 19007 0 1 3127
box 0 0 1 1
use contact_7  contact_7_119
timestamp 1634918361
transform 1 0 17839 0 1 3127
box 0 0 1 1
use contact_7  contact_7_120
timestamp 1634918361
transform 1 0 16671 0 1 3127
box 0 0 1 1
use contact_7  contact_7_121
timestamp 1634918361
transform 1 0 15503 0 1 3127
box 0 0 1 1
use contact_7  contact_7_122
timestamp 1634918361
transform 1 0 6074 0 1 3232
box 0 0 1 1
use contact_7  contact_7_123
timestamp 1634918361
transform 1 0 2853 0 1 4827
box 0 0 1 1
use contact_7  contact_7_124
timestamp 1634918361
transform 1 0 2853 0 1 3127
box 0 0 1 1
use cr_1  cr_1_0
timestamp 1634918361
transform 1 0 9694 0 1 6838
box 2040 -3614 15038 1462
use contact_7  contact_7_125
timestamp 1634918361
transform 1 0 33606 0 1 9768
box 0 0 1 1
use contact_19  contact_19_238
timestamp 1634918361
transform 1 0 33607 0 1 9773
box 0 0 1 1
use contact_7  contact_7_126
timestamp 1634918361
transform 1 0 34184 0 1 9768
box 0 0 1 1
use contact_7  contact_7_127
timestamp 1634918361
transform 1 0 33686 0 1 11326
box 0 0 1 1
use contact_19  contact_19_239
timestamp 1634918361
transform 1 0 33687 0 1 11331
box 0 0 1 1
use contact_7  contact_7_128
timestamp 1634918361
transform 1 0 34184 0 1 11326
box 0 0 1 1
use contact_7  contact_7_129
timestamp 1634918361
transform 1 0 33766 0 1 12596
box 0 0 1 1
use contact_19  contact_19_240
timestamp 1634918361
transform 1 0 33767 0 1 12601
box 0 0 1 1
use contact_7  contact_7_130
timestamp 1634918361
transform 1 0 34184 0 1 12596
box 0 0 1 1
use contact_7  contact_7_131
timestamp 1634918361
transform 1 0 33846 0 1 14154
box 0 0 1 1
use contact_19  contact_19_241
timestamp 1634918361
transform 1 0 33847 0 1 14159
box 0 0 1 1
use contact_7  contact_7_132
timestamp 1634918361
transform 1 0 34184 0 1 14154
box 0 0 1 1
use contact_7  contact_7_133
timestamp 1634918361
transform 1 0 9934 0 1 26126
box 0 0 1 1
use contact_19  contact_19_242
timestamp 1634918361
transform 1 0 9935 0 1 26131
box 0 0 1 1
use contact_7  contact_7_134
timestamp 1634918361
transform 1 0 9440 0 1 26126
box 0 0 1 1
use contact_7  contact_7_135
timestamp 1634918361
transform 1 0 9854 0 1 24568
box 0 0 1 1
use contact_19  contact_19_243
timestamp 1634918361
transform 1 0 9855 0 1 24573
box 0 0 1 1
use contact_7  contact_7_136
timestamp 1634918361
transform 1 0 9440 0 1 24568
box 0 0 1 1
use contact_7  contact_7_137
timestamp 1634918361
transform 1 0 9774 0 1 23298
box 0 0 1 1
use contact_19  contact_19_244
timestamp 1634918361
transform 1 0 9775 0 1 23303
box 0 0 1 1
use contact_7  contact_7_138
timestamp 1634918361
transform 1 0 9440 0 1 23298
box 0 0 1 1
use contact_7  contact_7_139
timestamp 1634918361
transform 1 0 9694 0 1 21740
box 0 0 1 1
use contact_19  contact_19_245
timestamp 1634918361
transform 1 0 9695 0 1 21745
box 0 0 1 1
use contact_7  contact_7_140
timestamp 1634918361
transform 1 0 9440 0 1 21740
box 0 0 1 1
use contact_30  contact_30_598
timestamp 1634918361
transform 1 0 40787 0 1 12798
box 0 0 1 1
use contact_7  contact_7_141
timestamp 1634918361
transform 1 0 40792 0 1 12794
box 0 0 1 1
use contact_30  contact_30_599
timestamp 1634918361
transform 1 0 40787 0 1 23033
box 0 0 1 1
use contact_30  contact_30_600
timestamp 1634918361
transform 1 0 2635 0 1 20280
box 0 0 1 1
use contact_7  contact_7_142
timestamp 1634918361
transform 1 0 2640 0 1 20276
box 0 0 1 1
use contact_30  contact_30_601
timestamp 1634918361
transform 1 0 2635 0 1 12873
box 0 0 1 1
use contact_7  contact_7_143
timestamp 1634918361
transform 1 0 27897 0 1 22730
box 0 0 1 1
use contact_7  contact_7_144
timestamp 1634918361
transform 1 0 34131 0 1 22730
box 0 0 1 1
use contact_7  contact_7_145
timestamp 1634918361
transform 1 0 26088 0 1 24181
box 0 0 1 1
use contact_7  contact_7_146
timestamp 1634918361
transform 1 0 34131 0 1 24181
box 0 0 1 1
use contact_7  contact_7_147
timestamp 1634918361
transform 1 0 25964 0 1 25542
box 0 0 1 1
use contact_7  contact_7_148
timestamp 1634918361
transform 1 0 34131 0 1 25542
box 0 0 1 1
use contact_7  contact_7_149
timestamp 1634918361
transform 1 0 15643 0 1 13168
box 0 0 1 1
use contact_7  contact_7_150
timestamp 1634918361
transform 1 0 9493 0 1 13168
box 0 0 1 1
use contact_7  contact_7_151
timestamp 1634918361
transform 1 0 17294 0 1 10377
box 0 0 1 1
use contact_7  contact_7_152
timestamp 1634918361
transform 1 0 9493 0 1 10377
box 0 0 1 1
use contact_7  contact_7_153
timestamp 1634918361
transform 1 0 17542 0 1 8926
box 0 0 1 1
use contact_7  contact_7_154
timestamp 1634918361
transform 1 0 9493 0 1 8926
box 0 0 1 1
use contact_7  contact_7_155
timestamp 1634918361
transform 1 0 17418 0 1 7528
box 0 0 1 1
use contact_7  contact_7_156
timestamp 1634918361
transform 1 0 9493 0 1 7528
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1634918361
transform 1 0 34047 0 1 14481
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1634918361
transform 1 0 9577 0 1 2871
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1634918361
transform 1 0 9577 0 1 21413
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1634918361
transform 1 0 15366 0 1 2600
box -36 -49 9380 1467
use wmask_dff  wmask_dff_0
timestamp 1634918361
transform 1 0 10694 0 1 2600
box -36 -49 4708 1467
use row_addr_dff  row_addr_dff_0
timestamp 1634918361
transform -1 0 35332 0 -1 14826
box -36 -49 1204 5705
use row_addr_dff  row_addr_dff_1
timestamp 1634918361
transform 1 0 8358 0 1 21142
box -36 -49 1204 5705
use control_logic_r  control_logic_r_0
timestamp 1634918361
transform -1 0 40782 0 -1 30544
box -75 -49 6618 18431
use control_logic_rw  control_logic_rw_0
timestamp 1634918361
transform 1 0 2716 0 1 2600
box -75 -49 6810 18431
use bank  bank_0
timestamp 1634918361
transform 1 0 9694 0 1 6838
box 0 0 24302 18696
<< labels >>
rlabel metal3 s 0 2992 212 3068 4 csb0
port 1 nsew
rlabel metal3 s 0 4760 212 4836 4 web0
port 2 nsew
rlabel metal4 s 5984 0 6060 212 4 clk0
port 3 nsew
rlabel metal4 s 15504 0 15580 212 4 din0[0]
port 4 nsew
rlabel metal4 s 16728 0 16804 212 4 din0[1]
port 5 nsew
rlabel metal4 s 17952 0 18028 212 4 din0[2]
port 6 nsew
rlabel metal4 s 19040 0 19116 212 4 din0[3]
port 7 nsew
rlabel metal4 s 20264 0 20340 212 4 din0[4]
port 8 nsew
rlabel metal4 s 21352 0 21428 212 4 din0[5]
port 9 nsew
rlabel metal4 s 22576 0 22652 212 4 din0[6]
port 10 nsew
rlabel metal4 s 23800 0 23876 212 4 din0[7]
port 11 nsew
rlabel metal4 s 19720 0 19796 212 4 dout0[0]
port 12 nsew
rlabel metal4 s 20400 0 20476 212 4 dout0[1]
port 13 nsew
rlabel metal4 s 20944 0 21020 212 4 dout0[2]
port 14 nsew
rlabel metal4 s 21624 0 21700 212 4 dout0[3]
port 15 nsew
rlabel metal4 s 22440 0 22516 212 4 dout0[4]
port 16 nsew
rlabel metal4 s 22848 0 22924 212 4 dout0[5]
port 17 nsew
rlabel metal4 s 23664 0 23740 212 4 dout0[6]
port 18 nsew
rlabel metal4 s 24072 0 24148 212 4 dout0[7]
port 19 nsew
rlabel metal3 s 0 21624 212 21700 4 addr0[0]
port 20 nsew
rlabel metal3 s 0 23256 212 23332 4 addr0[1]
port 21 nsew
rlabel metal3 s 0 24616 212 24692 4 addr0[2]
port 22 nsew
rlabel metal4 s 8568 32912 8644 33124 4 addr0[3]
port 23 nsew
rlabel metal4 s 10744 0 10820 212 4 wmask0[0]
port 24 nsew
rlabel metal4 s 12104 0 12180 212 4 wmask0[1]
port 25 nsew
rlabel metal4 s 13192 0 13268 212 4 wmask0[2]
port 26 nsew
rlabel metal4 s 14416 0 14492 212 4 wmask0[3]
port 27 nsew
rlabel metal3 s 43248 30056 43460 30132 4 csb1
port 28 nsew
rlabel metal4 s 37400 32912 37476 33124 4 clk1
port 29 nsew
rlabel metal4 s 19312 32912 19388 33124 4 dout1[0]
port 30 nsew
rlabel metal4 s 20400 32912 20476 33124 4 dout1[1]
port 31 nsew
rlabel metal4 s 20672 32912 20748 33124 4 dout1[2]
port 32 nsew
rlabel metal4 s 21624 32912 21700 33124 4 dout1[3]
port 33 nsew
rlabel metal4 s 21896 32912 21972 33124 4 dout1[4]
port 34 nsew
rlabel metal4 s 22848 32912 22924 33124 4 dout1[5]
port 35 nsew
rlabel metal4 s 23120 32912 23196 33124 4 dout1[6]
port 36 nsew
rlabel metal4 s 24208 32912 24284 33124 4 dout1[7]
port 37 nsew
rlabel metal3 s 43248 14144 43460 14220 4 addr1[0]
port 38 nsew
rlabel metal3 s 43248 12648 43460 12724 4 addr1[1]
port 39 nsew
rlabel metal3 s 43248 11288 43460 11364 4 addr1[2]
port 40 nsew
rlabel metal3 s 43248 9656 43460 9732 4 addr1[3]
port 41 nsew
rlabel metal3 s 952 952 42508 1300 4 vccd1
port 42 nsew
rlabel metal4 s 952 952 1300 32172 4 vccd1
port 42 nsew
rlabel metal4 s 42160 952 42508 32172 4 vccd1
port 42 nsew
rlabel metal3 s 952 31824 42508 32172 4 vccd1
port 42 nsew
rlabel metal3 s 272 272 43188 620 4 vssd1
port 43 nsew
rlabel metal4 s 42840 272 43188 32852 4 vssd1
port 43 nsew
rlabel metal3 s 272 32504 43188 32852 4 vssd1
port 43 nsew
rlabel metal4 s 272 272 620 32852 4 vssd1
port 43 nsew
<< properties >>
string FIXED_BBOX 0 0 43460 33124
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 362744
string GDS_START 132
<< end >>
