magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1309 -1260 9049 9160
<< metal1 >>
rect -32 7431 -26 7483
rect 26 7431 32 7483
rect -32 637 -26 689
rect 26 637 32 689
rect 972 0 1008 7900
rect 1044 0 1080 7900
rect 1116 7189 1152 7530
rect 1116 6399 1152 7031
rect 1116 5609 1152 6241
rect 1116 4819 1152 5451
rect 1116 4029 1152 4661
rect 1116 3239 1152 3871
rect 1116 2449 1152 3081
rect 1116 1659 1152 2291
rect 1116 869 1152 1501
rect 1116 370 1152 711
rect 1188 0 1224 7900
rect 1260 0 1296 7900
rect 1452 0 1488 7900
rect 1524 0 1560 7900
rect 1668 0 1704 7900
rect 1740 0 1776 7900
rect 2220 0 2256 7900
rect 2292 0 2328 7900
rect 2436 0 2472 7900
rect 2508 0 2544 7900
rect 2700 0 2736 7900
rect 2772 0 2808 7900
rect 2916 0 2952 7900
rect 2988 0 3024 7900
rect 3468 0 3504 7900
rect 3540 0 3576 7900
rect 3684 0 3720 7900
rect 3756 0 3792 7900
rect 3948 0 3984 7900
rect 4020 0 4056 7900
rect 4164 0 4200 7900
rect 4236 0 4272 7900
rect 4716 0 4752 7900
rect 4788 0 4824 7900
rect 4932 0 4968 7900
rect 5004 0 5040 7900
rect 5196 0 5232 7900
rect 5268 0 5304 7900
rect 5412 0 5448 7900
rect 5484 0 5520 7900
rect 5964 0 6000 7900
rect 6036 0 6072 7900
rect 6180 0 6216 7900
rect 6252 0 6288 7900
rect 6444 0 6480 7900
rect 6516 0 6552 7900
rect 6588 7189 6624 7530
rect 6588 6399 6624 7031
rect 6588 5609 6624 6241
rect 6588 4819 6624 5451
rect 6588 4029 6624 4661
rect 6588 3239 6624 3871
rect 6588 2449 6624 3081
rect 6588 1659 6624 2291
rect 6588 869 6624 1501
rect 6588 370 6624 711
rect 6660 0 6696 7900
rect 6732 0 6768 7900
rect 7708 7431 7714 7483
rect 7766 7431 7772 7483
rect 7708 637 7714 689
rect 7766 637 7772 689
<< via1 >>
rect -26 7431 26 7483
rect -26 637 26 689
rect 7714 7431 7766 7483
rect 7714 637 7766 689
<< metal2 >>
rect -37 7429 -28 7485
rect 28 7481 37 7485
rect 7703 7481 7712 7485
rect 28 7433 7712 7481
rect 28 7429 37 7433
rect 7703 7429 7712 7433
rect 7768 7429 7777 7485
rect 1080 7309 1188 7385
rect 6552 7309 6660 7385
rect 0 7213 7740 7261
rect 1080 7055 1188 7165
rect 6552 7055 6660 7165
rect 0 6959 7740 7007
rect 1080 6835 1188 6911
rect 6552 6835 6660 6911
rect 0 6739 7740 6787
rect 0 6643 7740 6691
rect 1080 6519 1188 6595
rect 6552 6519 6660 6595
rect 0 6423 7740 6471
rect 1080 6265 1188 6375
rect 6552 6265 6660 6375
rect 0 6169 7740 6217
rect 1080 6045 1188 6121
rect 6552 6045 6660 6121
rect 0 5949 7740 5997
rect 0 5853 7740 5901
rect 1080 5729 1188 5805
rect 6552 5729 6660 5805
rect 0 5633 7740 5681
rect 1080 5475 1188 5585
rect 6552 5475 6660 5585
rect 0 5379 7740 5427
rect 1080 5255 1188 5331
rect 6552 5255 6660 5331
rect 0 5159 7740 5207
rect 0 5063 7740 5111
rect 1080 4939 1188 5015
rect 6552 4939 6660 5015
rect 0 4843 7740 4891
rect 1080 4685 1188 4795
rect 6552 4685 6660 4795
rect 0 4589 7740 4637
rect 1080 4465 1188 4541
rect 6552 4465 6660 4541
rect 0 4369 7740 4417
rect 0 4273 7740 4321
rect 1080 4149 1188 4225
rect 6552 4149 6660 4225
rect 0 4053 7740 4101
rect 1080 3895 1188 4005
rect 6552 3895 6660 4005
rect 0 3799 7740 3847
rect 1080 3675 1188 3751
rect 6552 3675 6660 3751
rect 0 3579 7740 3627
rect 0 3483 7740 3531
rect 1080 3359 1188 3435
rect 6552 3359 6660 3435
rect 0 3263 7740 3311
rect 1080 3105 1188 3215
rect 6552 3105 6660 3215
rect 0 3009 7740 3057
rect 1080 2885 1188 2961
rect 6552 2885 6660 2961
rect 0 2789 7740 2837
rect 0 2693 7740 2741
rect 1080 2569 1188 2645
rect 6552 2569 6660 2645
rect 0 2473 7740 2521
rect 1080 2315 1188 2425
rect 6552 2315 6660 2425
rect 0 2219 7740 2267
rect 1080 2095 1188 2171
rect 6552 2095 6660 2171
rect 0 1999 7740 2047
rect 0 1903 7740 1951
rect 1080 1779 1188 1855
rect 6552 1779 6660 1855
rect 0 1683 7740 1731
rect 1080 1525 1188 1635
rect 6552 1525 6660 1635
rect 0 1429 7740 1477
rect 1080 1305 1188 1381
rect 6552 1305 6660 1381
rect 0 1209 7740 1257
rect 0 1113 7740 1161
rect 1080 989 1188 1065
rect 6552 989 6660 1065
rect 0 893 7740 941
rect 1080 735 1188 845
rect 6552 735 6660 845
rect -37 635 -28 691
rect 28 687 37 691
rect 7703 687 7712 691
rect 28 639 7712 687
rect 28 635 37 639
rect 7703 635 7712 639
rect 7768 635 7777 691
rect 1080 515 1188 591
rect 6552 515 6660 591
rect 0 419 7740 467
<< via2 >>
rect -28 7483 28 7485
rect -28 7431 -26 7483
rect -26 7431 26 7483
rect 26 7431 28 7483
rect 7712 7483 7768 7485
rect -28 7429 28 7431
rect 7712 7431 7714 7483
rect 7714 7431 7766 7483
rect 7766 7431 7768 7483
rect 7712 7429 7768 7431
rect -28 689 28 691
rect -28 637 -26 689
rect -26 637 26 689
rect 26 637 28 689
rect 7712 689 7768 691
rect -28 635 28 637
rect 7712 637 7714 689
rect 7714 637 7766 689
rect 7766 637 7768 689
rect 7712 635 7768 637
<< metal3 >>
rect 1013 7622 1111 7720
rect 1637 7622 1735 7720
rect 2261 7622 2359 7720
rect 2885 7622 2983 7720
rect 3509 7622 3607 7720
rect 4133 7622 4231 7720
rect 4757 7622 4855 7720
rect 5381 7622 5479 7720
rect 6005 7622 6103 7720
rect 6629 7622 6727 7720
rect -49 7485 49 7506
rect -49 7429 -28 7485
rect 28 7429 49 7485
rect -49 7408 49 7429
rect 7691 7485 7789 7506
rect 7691 7429 7712 7485
rect 7768 7429 7789 7485
rect 7691 7408 7789 7429
rect 317 7061 415 7159
rect 7325 7061 7423 7159
rect 317 6824 415 6922
rect 7325 6824 7423 6922
rect 317 6508 415 6606
rect 7325 6508 7423 6606
rect 317 6271 415 6369
rect 7325 6271 7423 6369
rect 317 6034 415 6132
rect 7325 6034 7423 6132
rect 317 5718 415 5816
rect 7325 5718 7423 5816
rect 317 5481 415 5579
rect 7325 5481 7423 5579
rect 317 5244 415 5342
rect 7325 5244 7423 5342
rect 317 4928 415 5026
rect 7325 4928 7423 5026
rect 317 4691 415 4789
rect 7325 4691 7423 4789
rect 317 4454 415 4552
rect 7325 4454 7423 4552
rect 317 4138 415 4236
rect 7325 4138 7423 4236
rect 317 3901 415 3999
rect 7325 3901 7423 3999
rect 317 3664 415 3762
rect 7325 3664 7423 3762
rect 317 3348 415 3446
rect 7325 3348 7423 3446
rect 317 3111 415 3209
rect 7325 3111 7423 3209
rect 317 2874 415 2972
rect 7325 2874 7423 2972
rect 317 2558 415 2656
rect 7325 2558 7423 2656
rect 317 2321 415 2419
rect 7325 2321 7423 2419
rect 317 2084 415 2182
rect 7325 2084 7423 2182
rect 317 1768 415 1866
rect 7325 1768 7423 1866
rect 317 1531 415 1629
rect 7325 1531 7423 1629
rect 317 1294 415 1392
rect 7325 1294 7423 1392
rect 317 978 415 1076
rect 7325 978 7423 1076
rect 317 741 415 839
rect 7325 741 7423 839
rect -49 691 49 712
rect -49 635 -28 691
rect 28 635 49 691
rect -49 614 49 635
rect 7691 691 7789 712
rect 7691 635 7712 691
rect 7768 635 7789 691
rect 7691 614 7789 635
rect 1013 180 1111 278
rect 1637 180 1735 278
rect 2261 180 2359 278
rect 2885 180 2983 278
rect 3509 180 3607 278
rect 4133 180 4231 278
rect 4757 180 4855 278
rect 5381 180 5479 278
rect 6005 180 6103 278
rect 6629 180 6727 278
use contact_9  contact_9_0
timestamp 1634918361
transform 1 0 7703 0 1 7424
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1634918361
transform 1 0 7708 0 1 7431
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1634918361
transform 1 0 -37 0 1 7424
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1634918361
transform 1 0 -32 0 1 7431
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1634918361
transform 1 0 7703 0 1 630
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1634918361
transform 1 0 7708 0 1 637
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1634918361
transform 1 0 -37 0 1 630
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1634918361
transform 1 0 -32 0 1 637
box 0 0 1 1
use row_cap_array_0  row_cap_array_0_0
timestamp 1634918361
transform 1 0 6990 0 1 0
box 0 419 666 7481
use row_cap_array  row_cap_array_0
timestamp 1634918361
transform 1 0 126 0 1 0
box -42 419 624 7481
use col_cap_array  col_cap_array_0
timestamp 1634918361
transform 1 0 1374 0 -1 7900
box 0 0 4992 474
use col_cap_array_0  col_cap_array_0_0
timestamp 1634918361
transform 1 0 1374 0 1 0
box 0 0 4992 474
use dummy_array  dummy_array_0
timestamp 1634918361
transform 1 0 1374 0 1 7110
box -42 -105 5034 421
use dummy_array  dummy_array_1
timestamp 1634918361
transform 1 0 1374 0 -1 790
box -42 -105 5034 421
use replica_column_0  replica_column_0_0
timestamp 1634918361
transform 1 0 6366 0 1 0
box -42 0 650 7900
use replica_column  replica_column_0
timestamp 1634918361
transform 1 0 750 0 1 0
box -26 0 666 7900
use bitcell_array  bitcell_array_0
timestamp 1634918361
transform 1 0 1374 0 1 790
box -42 -105 5034 6425
<< labels >>
rlabel metal2 s 0 1113 7740 1161 4 wl_0_0
port 1 nsew
rlabel metal2 s 0 893 7740 941 4 wl_1_0
port 2 nsew
rlabel metal2 s 0 1209 7740 1257 4 wl_0_1
port 3 nsew
rlabel metal2 s 0 1429 7740 1477 4 wl_1_1
port 4 nsew
rlabel metal2 s 0 1903 7740 1951 4 wl_0_2
port 5 nsew
rlabel metal2 s 0 1683 7740 1731 4 wl_1_2
port 6 nsew
rlabel metal2 s 0 1999 7740 2047 4 wl_0_3
port 7 nsew
rlabel metal2 s 0 2219 7740 2267 4 wl_1_3
port 8 nsew
rlabel metal2 s 0 2693 7740 2741 4 wl_0_4
port 9 nsew
rlabel metal2 s 0 2473 7740 2521 4 wl_1_4
port 10 nsew
rlabel metal2 s 0 2789 7740 2837 4 wl_0_5
port 11 nsew
rlabel metal2 s 0 3009 7740 3057 4 wl_1_5
port 12 nsew
rlabel metal2 s 0 3483 7740 3531 4 wl_0_6
port 13 nsew
rlabel metal2 s 0 3263 7740 3311 4 wl_1_6
port 14 nsew
rlabel metal2 s 0 3579 7740 3627 4 wl_0_7
port 15 nsew
rlabel metal2 s 0 3799 7740 3847 4 wl_1_7
port 16 nsew
rlabel metal2 s 0 4273 7740 4321 4 wl_0_8
port 17 nsew
rlabel metal2 s 0 4053 7740 4101 4 wl_1_8
port 18 nsew
rlabel metal2 s 0 4369 7740 4417 4 wl_0_9
port 19 nsew
rlabel metal2 s 0 4589 7740 4637 4 wl_1_9
port 20 nsew
rlabel metal2 s 0 5063 7740 5111 4 wl_0_10
port 21 nsew
rlabel metal2 s 0 4843 7740 4891 4 wl_1_10
port 22 nsew
rlabel metal2 s 0 5159 7740 5207 4 wl_0_11
port 23 nsew
rlabel metal2 s 0 5379 7740 5427 4 wl_1_11
port 24 nsew
rlabel metal2 s 0 5853 7740 5901 4 wl_0_12
port 25 nsew
rlabel metal2 s 0 5633 7740 5681 4 wl_1_12
port 26 nsew
rlabel metal2 s 0 5949 7740 5997 4 wl_0_13
port 27 nsew
rlabel metal2 s 0 6169 7740 6217 4 wl_1_13
port 28 nsew
rlabel metal2 s 0 6643 7740 6691 4 wl_0_14
port 29 nsew
rlabel metal2 s 0 6423 7740 6471 4 wl_1_14
port 30 nsew
rlabel metal2 s 0 6739 7740 6787 4 wl_0_15
port 31 nsew
rlabel metal2 s 0 6959 7740 7007 4 wl_1_15
port 32 nsew
rlabel metal2 s 0 419 7740 467 4 rbl_wl_0_0
port 33 nsew
rlabel metal2 s 0 7213 7740 7261 4 rbl_wl_1_1
port 34 nsew
rlabel metal1 s 1452 0 1488 7900 4 bl_0_0
port 35 nsew
rlabel metal1 s 1668 0 1704 7900 4 bl_1_0
port 36 nsew
rlabel metal1 s 1524 0 1560 7900 4 br_0_0
port 37 nsew
rlabel metal1 s 1740 0 1776 7900 4 br_1_0
port 38 nsew
rlabel metal1 s 2508 0 2544 7900 4 bl_0_1
port 39 nsew
rlabel metal1 s 2292 0 2328 7900 4 bl_1_1
port 40 nsew
rlabel metal1 s 2436 0 2472 7900 4 br_0_1
port 41 nsew
rlabel metal1 s 2220 0 2256 7900 4 br_1_1
port 42 nsew
rlabel metal1 s 2700 0 2736 7900 4 bl_0_2
port 43 nsew
rlabel metal1 s 2916 0 2952 7900 4 bl_1_2
port 44 nsew
rlabel metal1 s 2772 0 2808 7900 4 br_0_2
port 45 nsew
rlabel metal1 s 2988 0 3024 7900 4 br_1_2
port 46 nsew
rlabel metal1 s 3756 0 3792 7900 4 bl_0_3
port 47 nsew
rlabel metal1 s 3540 0 3576 7900 4 bl_1_3
port 48 nsew
rlabel metal1 s 3684 0 3720 7900 4 br_0_3
port 49 nsew
rlabel metal1 s 3468 0 3504 7900 4 br_1_3
port 50 nsew
rlabel metal1 s 3948 0 3984 7900 4 bl_0_4
port 51 nsew
rlabel metal1 s 4164 0 4200 7900 4 bl_1_4
port 52 nsew
rlabel metal1 s 4020 0 4056 7900 4 br_0_4
port 53 nsew
rlabel metal1 s 4236 0 4272 7900 4 br_1_4
port 54 nsew
rlabel metal1 s 5004 0 5040 7900 4 bl_0_5
port 55 nsew
rlabel metal1 s 4788 0 4824 7900 4 bl_1_5
port 56 nsew
rlabel metal1 s 4932 0 4968 7900 4 br_0_5
port 57 nsew
rlabel metal1 s 4716 0 4752 7900 4 br_1_5
port 58 nsew
rlabel metal1 s 5196 0 5232 7900 4 bl_0_6
port 59 nsew
rlabel metal1 s 5412 0 5448 7900 4 bl_1_6
port 60 nsew
rlabel metal1 s 5268 0 5304 7900 4 br_0_6
port 61 nsew
rlabel metal1 s 5484 0 5520 7900 4 br_1_6
port 62 nsew
rlabel metal1 s 6252 0 6288 7900 4 bl_0_7
port 63 nsew
rlabel metal1 s 6036 0 6072 7900 4 bl_1_7
port 64 nsew
rlabel metal1 s 6180 0 6216 7900 4 br_0_7
port 65 nsew
rlabel metal1 s 5964 0 6000 7900 4 br_1_7
port 66 nsew
rlabel metal1 s 1260 0 1296 7900 4 rbl_bl_0_0
port 67 nsew
rlabel metal1 s 1044 0 1080 7900 4 rbl_bl_1_0
port 68 nsew
rlabel metal1 s 1188 0 1224 7900 4 rbl_br_0_0
port 69 nsew
rlabel metal1 s 972 0 1008 7900 4 rbl_br_1_0
port 70 nsew
rlabel metal1 s 6444 0 6480 7900 4 rbl_bl_0_1
port 71 nsew
rlabel metal1 s 6660 0 6696 7900 4 rbl_bl_1_1
port 72 nsew
rlabel metal1 s 6516 0 6552 7900 4 rbl_br_0_1
port 73 nsew
rlabel metal1 s 6732 0 6768 7900 4 rbl_br_1_1
port 74 nsew
rlabel metal1 s 1116 7189 1152 7530 4 vdd
port 75 nsew
rlabel metal1 s 1116 1659 1152 2000 4 vdd
port 75 nsew
rlabel metal1 s 6588 2449 6624 2790 4 vdd
port 75 nsew
rlabel metal3 s 1013 180 1111 278 4 vdd
port 75 nsew
rlabel metal1 s 1116 4029 1152 4370 4 vdd
port 75 nsew
rlabel metal1 s 6588 6399 6624 6740 4 vdd
port 75 nsew
rlabel metal1 s 1116 4320 1152 4661 4 vdd
port 75 nsew
rlabel metal3 s 4133 7622 4231 7720 4 vdd
port 75 nsew
rlabel metal1 s 6588 869 6624 1210 4 vdd
port 75 nsew
rlabel metal1 s 6588 2740 6624 3081 4 vdd
port 75 nsew
rlabel metal3 s 3509 7622 3607 7720 4 vdd
port 75 nsew
rlabel metal1 s 6588 4029 6624 4370 4 vdd
port 75 nsew
rlabel metal3 s 5381 7622 5479 7720 4 vdd
port 75 nsew
rlabel metal1 s 6588 1950 6624 2291 4 vdd
port 75 nsew
rlabel metal1 s 6588 5609 6624 5950 4 vdd
port 75 nsew
rlabel metal1 s 1116 5609 1152 5950 4 vdd
port 75 nsew
rlabel metal1 s 1116 5900 1152 6241 4 vdd
port 75 nsew
rlabel metal1 s 6588 3530 6624 3871 4 vdd
port 75 nsew
rlabel metal3 s 1637 180 1735 278 4 vdd
port 75 nsew
rlabel metal3 s 2885 180 2983 278 4 vdd
port 75 nsew
rlabel metal3 s 2261 7622 2359 7720 4 vdd
port 75 nsew
rlabel metal1 s 1116 2449 1152 2790 4 vdd
port 75 nsew
rlabel metal1 s 6588 5110 6624 5451 4 vdd
port 75 nsew
rlabel metal1 s 6588 5900 6624 6241 4 vdd
port 75 nsew
rlabel metal1 s 6588 4320 6624 4661 4 vdd
port 75 nsew
rlabel metal3 s 6629 180 6727 278 4 vdd
port 75 nsew
rlabel metal1 s 6588 6690 6624 7031 4 vdd
port 75 nsew
rlabel metal1 s 6588 3239 6624 3580 4 vdd
port 75 nsew
rlabel metal3 s 3509 180 3607 278 4 vdd
port 75 nsew
rlabel metal3 s 1637 7622 1735 7720 4 vdd
port 75 nsew
rlabel metal3 s 6629 7622 6727 7720 4 vdd
port 75 nsew
rlabel metal1 s 6588 1659 6624 2000 4 vdd
port 75 nsew
rlabel metal3 s 4757 7622 4855 7720 4 vdd
port 75 nsew
rlabel metal3 s 6005 180 6103 278 4 vdd
port 75 nsew
rlabel metal3 s 6005 7622 6103 7720 4 vdd
port 75 nsew
rlabel metal1 s 1116 6399 1152 6740 4 vdd
port 75 nsew
rlabel metal1 s 6588 1160 6624 1501 4 vdd
port 75 nsew
rlabel metal1 s 6588 370 6624 711 4 vdd
port 75 nsew
rlabel metal3 s 5381 180 5479 278 4 vdd
port 75 nsew
rlabel metal3 s 2261 180 2359 278 4 vdd
port 75 nsew
rlabel metal1 s 1116 4819 1152 5160 4 vdd
port 75 nsew
rlabel metal1 s 1116 1950 1152 2291 4 vdd
port 75 nsew
rlabel metal1 s 1116 2740 1152 3081 4 vdd
port 75 nsew
rlabel metal1 s 1116 3239 1152 3580 4 vdd
port 75 nsew
rlabel metal3 s 4757 180 4855 278 4 vdd
port 75 nsew
rlabel metal1 s 1116 370 1152 711 4 vdd
port 75 nsew
rlabel metal1 s 6588 4819 6624 5160 4 vdd
port 75 nsew
rlabel metal1 s 1116 3530 1152 3871 4 vdd
port 75 nsew
rlabel metal1 s 1116 6690 1152 7031 4 vdd
port 75 nsew
rlabel metal3 s 2885 7622 2983 7720 4 vdd
port 75 nsew
rlabel metal1 s 6588 7189 6624 7530 4 vdd
port 75 nsew
rlabel metal3 s 4133 180 4231 278 4 vdd
port 75 nsew
rlabel metal1 s 1116 1160 1152 1501 4 vdd
port 75 nsew
rlabel metal1 s 1116 869 1152 1210 4 vdd
port 75 nsew
rlabel metal3 s 1013 7622 1111 7720 4 vdd
port 75 nsew
rlabel metal1 s 1116 5110 1152 5451 4 vdd
port 75 nsew
rlabel metal2 s 1080 2315 1188 2425 4 gnd
port 76 nsew
rlabel metal3 s 7325 2084 7423 2182 4 gnd
port 76 nsew
rlabel metal3 s 317 3664 415 3762 4 gnd
port 76 nsew
rlabel metal3 s 7325 1294 7423 1392 4 gnd
port 76 nsew
rlabel metal2 s 1080 4465 1188 4541 4 gnd
port 76 nsew
rlabel metal3 s 317 1294 415 1392 4 gnd
port 76 nsew
rlabel metal2 s 1080 1525 1188 1635 4 gnd
port 76 nsew
rlabel metal3 s 7325 1531 7423 1629 4 gnd
port 76 nsew
rlabel metal2 s 6552 6045 6660 6121 4 gnd
port 76 nsew
rlabel metal3 s 7325 2321 7423 2419 4 gnd
port 76 nsew
rlabel metal3 s 7325 978 7423 1076 4 gnd
port 76 nsew
rlabel metal3 s 317 1768 415 1866 4 gnd
port 76 nsew
rlabel metal3 s 7325 1768 7423 1866 4 gnd
port 76 nsew
rlabel metal2 s 6552 6835 6660 6911 4 gnd
port 76 nsew
rlabel metal3 s 7325 5718 7423 5816 4 gnd
port 76 nsew
rlabel metal2 s 6552 5255 6660 5331 4 gnd
port 76 nsew
rlabel metal2 s 1080 3359 1188 3435 4 gnd
port 76 nsew
rlabel metal2 s 6552 6519 6660 6595 4 gnd
port 76 nsew
rlabel metal3 s -49 614 49 712 4 gnd
port 76 nsew
rlabel metal2 s 1080 5475 1188 5585 4 gnd
port 76 nsew
rlabel metal3 s 7325 3111 7423 3209 4 gnd
port 76 nsew
rlabel metal2 s 1080 3105 1188 3215 4 gnd
port 76 nsew
rlabel metal2 s 1080 7055 1188 7165 4 gnd
port 76 nsew
rlabel metal2 s 6552 7309 6660 7385 4 gnd
port 76 nsew
rlabel metal2 s 1080 5729 1188 5805 4 gnd
port 76 nsew
rlabel metal2 s 1080 989 1188 1065 4 gnd
port 76 nsew
rlabel metal3 s 7325 4138 7423 4236 4 gnd
port 76 nsew
rlabel metal2 s 1080 4939 1188 5015 4 gnd
port 76 nsew
rlabel metal3 s 317 7061 415 7159 4 gnd
port 76 nsew
rlabel metal3 s 317 978 415 1076 4 gnd
port 76 nsew
rlabel metal3 s 7325 4928 7423 5026 4 gnd
port 76 nsew
rlabel metal3 s 7325 3664 7423 3762 4 gnd
port 76 nsew
rlabel metal3 s 317 6824 415 6922 4 gnd
port 76 nsew
rlabel metal2 s 1080 6519 1188 6595 4 gnd
port 76 nsew
rlabel metal3 s 317 741 415 839 4 gnd
port 76 nsew
rlabel metal2 s 6552 1779 6660 1855 4 gnd
port 76 nsew
rlabel metal3 s 7325 7061 7423 7159 4 gnd
port 76 nsew
rlabel metal2 s 6552 4685 6660 4795 4 gnd
port 76 nsew
rlabel metal2 s 1080 5255 1188 5331 4 gnd
port 76 nsew
rlabel metal2 s 1080 515 1188 591 4 gnd
port 76 nsew
rlabel metal3 s 7691 614 7789 712 4 gnd
port 76 nsew
rlabel metal2 s 1080 6045 1188 6121 4 gnd
port 76 nsew
rlabel metal3 s 7325 4691 7423 4789 4 gnd
port 76 nsew
rlabel metal2 s 1080 7309 1188 7385 4 gnd
port 76 nsew
rlabel metal3 s 317 4454 415 4552 4 gnd
port 76 nsew
rlabel metal2 s 1080 6835 1188 6911 4 gnd
port 76 nsew
rlabel metal3 s -49 7408 49 7506 4 gnd
port 76 nsew
rlabel metal3 s 317 2558 415 2656 4 gnd
port 76 nsew
rlabel metal2 s 6552 3359 6660 3435 4 gnd
port 76 nsew
rlabel metal2 s 6552 3105 6660 3215 4 gnd
port 76 nsew
rlabel metal3 s 317 5718 415 5816 4 gnd
port 76 nsew
rlabel metal3 s 317 6271 415 6369 4 gnd
port 76 nsew
rlabel metal3 s 7325 6508 7423 6606 4 gnd
port 76 nsew
rlabel metal2 s 1080 6265 1188 6375 4 gnd
port 76 nsew
rlabel metal3 s 317 5244 415 5342 4 gnd
port 76 nsew
rlabel metal3 s 7325 3348 7423 3446 4 gnd
port 76 nsew
rlabel metal3 s 7325 6271 7423 6369 4 gnd
port 76 nsew
rlabel metal3 s 7691 7408 7789 7506 4 gnd
port 76 nsew
rlabel metal3 s 7325 5244 7423 5342 4 gnd
port 76 nsew
rlabel metal3 s 7325 2558 7423 2656 4 gnd
port 76 nsew
rlabel metal3 s 317 3348 415 3446 4 gnd
port 76 nsew
rlabel metal2 s 1080 2569 1188 2645 4 gnd
port 76 nsew
rlabel metal2 s 6552 515 6660 591 4 gnd
port 76 nsew
rlabel metal2 s 6552 3675 6660 3751 4 gnd
port 76 nsew
rlabel metal3 s 317 6034 415 6132 4 gnd
port 76 nsew
rlabel metal2 s 6552 2315 6660 2425 4 gnd
port 76 nsew
rlabel metal2 s 1080 3895 1188 4005 4 gnd
port 76 nsew
rlabel metal3 s 317 1531 415 1629 4 gnd
port 76 nsew
rlabel metal2 s 6552 6265 6660 6375 4 gnd
port 76 nsew
rlabel metal3 s 317 4691 415 4789 4 gnd
port 76 nsew
rlabel metal2 s 6552 3895 6660 4005 4 gnd
port 76 nsew
rlabel metal2 s 1080 3675 1188 3751 4 gnd
port 76 nsew
rlabel metal3 s 7325 6824 7423 6922 4 gnd
port 76 nsew
rlabel metal2 s 6552 4149 6660 4225 4 gnd
port 76 nsew
rlabel metal2 s 6552 989 6660 1065 4 gnd
port 76 nsew
rlabel metal2 s 6552 2569 6660 2645 4 gnd
port 76 nsew
rlabel metal3 s 317 6508 415 6606 4 gnd
port 76 nsew
rlabel metal2 s 6552 1305 6660 1381 4 gnd
port 76 nsew
rlabel metal3 s 7325 5481 7423 5579 4 gnd
port 76 nsew
rlabel metal2 s 6552 1525 6660 1635 4 gnd
port 76 nsew
rlabel metal3 s 317 4928 415 5026 4 gnd
port 76 nsew
rlabel metal2 s 6552 735 6660 845 4 gnd
port 76 nsew
rlabel metal2 s 6552 7055 6660 7165 4 gnd
port 76 nsew
rlabel metal2 s 1080 2885 1188 2961 4 gnd
port 76 nsew
rlabel metal3 s 317 3111 415 3209 4 gnd
port 76 nsew
rlabel metal3 s 317 5481 415 5579 4 gnd
port 76 nsew
rlabel metal2 s 1080 1305 1188 1381 4 gnd
port 76 nsew
rlabel metal3 s 7325 4454 7423 4552 4 gnd
port 76 nsew
rlabel metal2 s 6552 4465 6660 4541 4 gnd
port 76 nsew
rlabel metal3 s 317 2084 415 2182 4 gnd
port 76 nsew
rlabel metal3 s 317 4138 415 4236 4 gnd
port 76 nsew
rlabel metal2 s 1080 735 1188 845 4 gnd
port 76 nsew
rlabel metal3 s 7325 2874 7423 2972 4 gnd
port 76 nsew
rlabel metal3 s 317 3901 415 3999 4 gnd
port 76 nsew
rlabel metal2 s 6552 5475 6660 5585 4 gnd
port 76 nsew
rlabel metal2 s 1080 1779 1188 1855 4 gnd
port 76 nsew
rlabel metal3 s 7325 741 7423 839 4 gnd
port 76 nsew
rlabel metal2 s 6552 2885 6660 2961 4 gnd
port 76 nsew
rlabel metal2 s 6552 5729 6660 5805 4 gnd
port 76 nsew
rlabel metal3 s 7325 3901 7423 3999 4 gnd
port 76 nsew
rlabel metal2 s 1080 2095 1188 2171 4 gnd
port 76 nsew
rlabel metal2 s 6552 4939 6660 5015 4 gnd
port 76 nsew
rlabel metal3 s 317 2874 415 2972 4 gnd
port 76 nsew
rlabel metal2 s 6552 2095 6660 2171 4 gnd
port 76 nsew
rlabel metal2 s 1080 4149 1188 4225 4 gnd
port 76 nsew
rlabel metal3 s 317 2321 415 2419 4 gnd
port 76 nsew
rlabel metal3 s 7325 6034 7423 6132 4 gnd
port 76 nsew
rlabel metal2 s 1080 4685 1188 4795 4 gnd
port 76 nsew
<< properties >>
string FIXED_BBOX 0 0 7740 630
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 505204
string GDS_START 462346
<< end >>
