magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect 780 -4874 16298 2722
<< metal1 >>
rect 9866 1399 9872 1451
rect 9924 1399 9930 1451
rect 10420 1399 10426 1451
rect 10478 1399 10484 1451
rect 11114 1399 11120 1451
rect 11172 1399 11178 1451
rect 11668 1399 11674 1451
rect 11726 1399 11732 1451
rect 12362 1399 12368 1451
rect 12420 1399 12426 1451
rect 12916 1399 12922 1451
rect 12974 1399 12980 1451
rect 13610 1399 13616 1451
rect 13668 1399 13674 1451
rect 14164 1399 14170 1451
rect 14222 1399 14228 1451
<< via1 >>
rect 9872 1399 9924 1451
rect 10426 1399 10478 1451
rect 11120 1399 11172 1451
rect 11674 1399 11726 1451
rect 12368 1399 12420 1451
rect 12922 1399 12974 1451
rect 13616 1399 13668 1451
rect 14170 1399 14222 1451
<< metal2 >>
rect 9870 1453 9926 1462
rect 9870 1388 9926 1397
rect 10424 1453 10480 1462
rect 10424 1388 10480 1397
rect 11118 1453 11174 1462
rect 11118 1388 11174 1397
rect 11672 1453 11728 1462
rect 11672 1388 11728 1397
rect 12366 1453 12422 1462
rect 12366 1388 12422 1397
rect 12920 1453 12976 1462
rect 12920 1388 12976 1397
rect 13614 1453 13670 1462
rect 13614 1388 13670 1397
rect 14168 1453 14224 1462
rect 14168 1388 14224 1397
rect 9585 333 9641 342
rect 9585 268 9641 277
rect 10833 333 10889 342
rect 10833 268 10889 277
rect 12081 333 12137 342
rect 12081 268 12137 277
rect 13329 333 13385 342
rect 13329 268 13385 277
rect 2087 -3549 2143 -3540
rect 2087 -3614 2143 -3605
rect 3255 -3549 3311 -3540
rect 3255 -3614 3311 -3605
rect 4423 -3549 4479 -3540
rect 4423 -3614 4479 -3605
rect 5591 -3549 5647 -3540
rect 5591 -3614 5647 -3605
rect 6759 -3549 6815 -3540
rect 6759 -3614 6815 -3605
rect 7927 -3549 7983 -3540
rect 7927 -3614 7983 -3605
rect 9095 -3549 9151 -3540
rect 9095 -3614 9151 -3605
rect 10263 -3549 10319 -3540
rect 10263 -3614 10319 -3605
rect 11431 -3549 11487 -3540
rect 11431 -3614 11487 -3605
rect 12599 -3549 12655 -3540
rect 12599 -3614 12655 -3605
rect 13767 -3549 13823 -3540
rect 13767 -3614 13823 -3605
rect 14935 -3549 14991 -3540
rect 14935 -3614 14991 -3605
<< via2 >>
rect 9870 1451 9926 1453
rect 9870 1399 9872 1451
rect 9872 1399 9924 1451
rect 9924 1399 9926 1451
rect 9870 1397 9926 1399
rect 10424 1451 10480 1453
rect 10424 1399 10426 1451
rect 10426 1399 10478 1451
rect 10478 1399 10480 1451
rect 10424 1397 10480 1399
rect 11118 1451 11174 1453
rect 11118 1399 11120 1451
rect 11120 1399 11172 1451
rect 11172 1399 11174 1451
rect 11118 1397 11174 1399
rect 11672 1451 11728 1453
rect 11672 1399 11674 1451
rect 11674 1399 11726 1451
rect 11726 1399 11728 1451
rect 11672 1397 11728 1399
rect 12366 1451 12422 1453
rect 12366 1399 12368 1451
rect 12368 1399 12420 1451
rect 12420 1399 12422 1451
rect 12366 1397 12422 1399
rect 12920 1451 12976 1453
rect 12920 1399 12922 1451
rect 12922 1399 12974 1451
rect 12974 1399 12976 1451
rect 12920 1397 12976 1399
rect 13614 1451 13670 1453
rect 13614 1399 13616 1451
rect 13616 1399 13668 1451
rect 13668 1399 13670 1451
rect 13614 1397 13670 1399
rect 14168 1451 14224 1453
rect 14168 1399 14170 1451
rect 14170 1399 14222 1451
rect 14222 1399 14224 1451
rect 14168 1397 14224 1399
rect 9585 277 9641 333
rect 10833 277 10889 333
rect 12081 277 12137 333
rect 13329 277 13385 333
rect 2087 -3605 2143 -3549
rect 3255 -3605 3311 -3549
rect 4423 -3605 4479 -3549
rect 5591 -3605 5647 -3549
rect 6759 -3605 6815 -3549
rect 7927 -3605 7983 -3549
rect 9095 -3605 9151 -3549
rect 10263 -3605 10319 -3549
rect 11431 -3605 11487 -3549
rect 12599 -3605 12655 -3549
rect 13767 -3605 13823 -3549
rect 14935 -3605 14991 -3549
<< metal3 >>
rect 9865 1457 9931 1458
rect 10419 1457 10485 1458
rect 11113 1457 11179 1458
rect 11667 1457 11733 1458
rect 12361 1457 12427 1458
rect 12915 1457 12981 1458
rect 13609 1457 13675 1458
rect 14163 1457 14229 1458
rect 9823 1393 9866 1457
rect 9930 1393 9973 1457
rect 10377 1393 10420 1457
rect 10484 1393 10527 1457
rect 11071 1393 11114 1457
rect 11178 1393 11221 1457
rect 11625 1393 11668 1457
rect 11732 1393 11775 1457
rect 12319 1393 12362 1457
rect 12426 1393 12469 1457
rect 12873 1393 12916 1457
rect 12980 1393 13023 1457
rect 13567 1393 13610 1457
rect 13674 1393 13717 1457
rect 14121 1393 14164 1457
rect 14228 1393 14271 1457
rect 9865 1392 9931 1393
rect 10419 1392 10485 1393
rect 11113 1392 11179 1393
rect 11667 1392 11733 1393
rect 12361 1392 12427 1393
rect 12915 1392 12981 1393
rect 13609 1392 13675 1393
rect 14163 1392 14229 1393
rect 9580 337 9646 338
rect 10828 337 10894 338
rect 12076 337 12142 338
rect 13324 337 13390 338
rect 9538 273 9581 337
rect 9645 273 9688 337
rect 10786 273 10829 337
rect 10893 273 10936 337
rect 12034 273 12077 337
rect 12141 273 12184 337
rect 13282 273 13325 337
rect 13389 273 13432 337
rect 9580 272 9646 273
rect 10828 272 10894 273
rect 12076 272 12142 273
rect 13324 272 13390 273
rect 9085 -516 9091 -452
rect 9155 -454 9161 -452
rect 11108 -454 11114 -452
rect 9155 -514 11114 -454
rect 9155 -516 9161 -514
rect 11108 -516 11114 -514
rect 11178 -516 11184 -452
rect 7917 -760 7923 -696
rect 7987 -698 7993 -696
rect 10414 -698 10420 -696
rect 7987 -758 10420 -698
rect 7987 -760 7993 -758
rect 10414 -760 10420 -758
rect 10484 -760 10490 -696
rect 6749 -1004 6755 -940
rect 6819 -942 6825 -940
rect 9860 -942 9866 -940
rect 6819 -1002 9866 -942
rect 6819 -1004 6825 -1002
rect 9860 -1004 9866 -1002
rect 9930 -1004 9936 -940
rect 10253 -1004 10259 -940
rect 10323 -942 10329 -940
rect 11662 -942 11668 -940
rect 10323 -1002 11668 -942
rect 10323 -1004 10329 -1002
rect 11662 -1004 11668 -1002
rect 11732 -1004 11738 -940
rect 5581 -1248 5587 -1184
rect 5651 -1186 5657 -1184
rect 13319 -1186 13325 -1184
rect 5651 -1246 13325 -1186
rect 5651 -1248 5657 -1246
rect 13319 -1248 13325 -1246
rect 13389 -1248 13395 -1184
rect 4413 -1492 4419 -1428
rect 4483 -1430 4489 -1428
rect 12071 -1430 12077 -1428
rect 4483 -1490 12077 -1430
rect 4483 -1492 4489 -1490
rect 12071 -1492 12077 -1490
rect 12141 -1492 12147 -1428
rect 3245 -1736 3251 -1672
rect 3315 -1674 3321 -1672
rect 10823 -1674 10829 -1672
rect 3315 -1734 10829 -1674
rect 3315 -1736 3321 -1734
rect 10823 -1736 10829 -1734
rect 10893 -1736 10899 -1672
rect 11421 -1736 11427 -1672
rect 11491 -1674 11497 -1672
rect 12356 -1674 12362 -1672
rect 11491 -1734 12362 -1674
rect 11491 -1736 11497 -1734
rect 12356 -1736 12362 -1734
rect 12426 -1736 12432 -1672
rect 2077 -1980 2083 -1916
rect 2147 -1918 2153 -1916
rect 9575 -1918 9581 -1916
rect 2147 -1978 9581 -1918
rect 2147 -1980 2153 -1978
rect 9575 -1980 9581 -1978
rect 9645 -1980 9651 -1916
rect 12589 -1980 12595 -1916
rect 12659 -1918 12665 -1916
rect 12910 -1918 12916 -1916
rect 12659 -1978 12916 -1918
rect 12659 -1980 12665 -1978
rect 12910 -1980 12916 -1978
rect 12980 -1980 12986 -1916
rect 13604 -1980 13610 -1916
rect 13674 -1918 13680 -1916
rect 13757 -1918 13763 -1916
rect 13674 -1978 13763 -1918
rect 13674 -1980 13680 -1978
rect 13757 -1980 13763 -1978
rect 13827 -1980 13833 -1916
rect 14158 -1980 14164 -1916
rect 14228 -1918 14234 -1916
rect 14925 -1918 14931 -1916
rect 14228 -1978 14931 -1918
rect 14228 -1980 14234 -1978
rect 14925 -1980 14931 -1978
rect 14995 -1980 15001 -1916
rect 2082 -3545 2148 -3544
rect 3250 -3545 3316 -3544
rect 4418 -3545 4484 -3544
rect 5586 -3545 5652 -3544
rect 6754 -3545 6820 -3544
rect 7922 -3545 7988 -3544
rect 9090 -3545 9156 -3544
rect 10258 -3545 10324 -3544
rect 11426 -3545 11492 -3544
rect 12594 -3545 12660 -3544
rect 13762 -3545 13828 -3544
rect 14930 -3545 14996 -3544
rect 2040 -3609 2083 -3545
rect 2147 -3609 2190 -3545
rect 3208 -3609 3251 -3545
rect 3315 -3609 3358 -3545
rect 4376 -3609 4419 -3545
rect 4483 -3609 4526 -3545
rect 5544 -3609 5587 -3545
rect 5651 -3609 5694 -3545
rect 6712 -3609 6755 -3545
rect 6819 -3609 6862 -3545
rect 7880 -3609 7923 -3545
rect 7987 -3609 8030 -3545
rect 9048 -3609 9091 -3545
rect 9155 -3609 9198 -3545
rect 10216 -3609 10259 -3545
rect 10323 -3609 10366 -3545
rect 11384 -3609 11427 -3545
rect 11491 -3609 11534 -3545
rect 12552 -3609 12595 -3545
rect 12659 -3609 12702 -3545
rect 13720 -3609 13763 -3545
rect 13827 -3609 13870 -3545
rect 14888 -3609 14931 -3545
rect 14995 -3609 15038 -3545
rect 2082 -3610 2148 -3609
rect 3250 -3610 3316 -3609
rect 4418 -3610 4484 -3609
rect 5586 -3610 5652 -3609
rect 6754 -3610 6820 -3609
rect 7922 -3610 7988 -3609
rect 9090 -3610 9156 -3609
rect 10258 -3610 10324 -3609
rect 11426 -3610 11492 -3609
rect 12594 -3610 12660 -3609
rect 13762 -3610 13828 -3609
rect 14930 -3610 14996 -3609
<< via3 >>
rect 9866 1453 9930 1457
rect 9866 1397 9870 1453
rect 9870 1397 9926 1453
rect 9926 1397 9930 1453
rect 9866 1393 9930 1397
rect 10420 1453 10484 1457
rect 10420 1397 10424 1453
rect 10424 1397 10480 1453
rect 10480 1397 10484 1453
rect 10420 1393 10484 1397
rect 11114 1453 11178 1457
rect 11114 1397 11118 1453
rect 11118 1397 11174 1453
rect 11174 1397 11178 1453
rect 11114 1393 11178 1397
rect 11668 1453 11732 1457
rect 11668 1397 11672 1453
rect 11672 1397 11728 1453
rect 11728 1397 11732 1453
rect 11668 1393 11732 1397
rect 12362 1453 12426 1457
rect 12362 1397 12366 1453
rect 12366 1397 12422 1453
rect 12422 1397 12426 1453
rect 12362 1393 12426 1397
rect 12916 1453 12980 1457
rect 12916 1397 12920 1453
rect 12920 1397 12976 1453
rect 12976 1397 12980 1453
rect 12916 1393 12980 1397
rect 13610 1453 13674 1457
rect 13610 1397 13614 1453
rect 13614 1397 13670 1453
rect 13670 1397 13674 1453
rect 13610 1393 13674 1397
rect 14164 1453 14228 1457
rect 14164 1397 14168 1453
rect 14168 1397 14224 1453
rect 14224 1397 14228 1453
rect 14164 1393 14228 1397
rect 9581 333 9645 337
rect 9581 277 9585 333
rect 9585 277 9641 333
rect 9641 277 9645 333
rect 9581 273 9645 277
rect 10829 333 10893 337
rect 10829 277 10833 333
rect 10833 277 10889 333
rect 10889 277 10893 333
rect 10829 273 10893 277
rect 12077 333 12141 337
rect 12077 277 12081 333
rect 12081 277 12137 333
rect 12137 277 12141 333
rect 12077 273 12141 277
rect 13325 333 13389 337
rect 13325 277 13329 333
rect 13329 277 13385 333
rect 13385 277 13389 333
rect 13325 273 13389 277
rect 9091 -516 9155 -452
rect 11114 -516 11178 -452
rect 7923 -760 7987 -696
rect 10420 -760 10484 -696
rect 6755 -1004 6819 -940
rect 9866 -1004 9930 -940
rect 10259 -1004 10323 -940
rect 11668 -1004 11732 -940
rect 5587 -1248 5651 -1184
rect 13325 -1248 13389 -1184
rect 4419 -1492 4483 -1428
rect 12077 -1492 12141 -1428
rect 3251 -1736 3315 -1672
rect 10829 -1736 10893 -1672
rect 11427 -1736 11491 -1672
rect 12362 -1736 12426 -1672
rect 2083 -1980 2147 -1916
rect 9581 -1980 9645 -1916
rect 12595 -1980 12659 -1916
rect 12916 -1980 12980 -1916
rect 13610 -1980 13674 -1916
rect 13763 -1980 13827 -1916
rect 14164 -1980 14228 -1916
rect 14931 -1980 14995 -1916
rect 2083 -3549 2147 -3545
rect 2083 -3605 2087 -3549
rect 2087 -3605 2143 -3549
rect 2143 -3605 2147 -3549
rect 2083 -3609 2147 -3605
rect 3251 -3549 3315 -3545
rect 3251 -3605 3255 -3549
rect 3255 -3605 3311 -3549
rect 3311 -3605 3315 -3549
rect 3251 -3609 3315 -3605
rect 4419 -3549 4483 -3545
rect 4419 -3605 4423 -3549
rect 4423 -3605 4479 -3549
rect 4479 -3605 4483 -3549
rect 4419 -3609 4483 -3605
rect 5587 -3549 5651 -3545
rect 5587 -3605 5591 -3549
rect 5591 -3605 5647 -3549
rect 5647 -3605 5651 -3549
rect 5587 -3609 5651 -3605
rect 6755 -3549 6819 -3545
rect 6755 -3605 6759 -3549
rect 6759 -3605 6815 -3549
rect 6815 -3605 6819 -3549
rect 6755 -3609 6819 -3605
rect 7923 -3549 7987 -3545
rect 7923 -3605 7927 -3549
rect 7927 -3605 7983 -3549
rect 7983 -3605 7987 -3549
rect 7923 -3609 7987 -3605
rect 9091 -3549 9155 -3545
rect 9091 -3605 9095 -3549
rect 9095 -3605 9151 -3549
rect 9151 -3605 9155 -3549
rect 9091 -3609 9155 -3605
rect 10259 -3549 10323 -3545
rect 10259 -3605 10263 -3549
rect 10263 -3605 10319 -3549
rect 10319 -3605 10323 -3549
rect 10259 -3609 10323 -3605
rect 11427 -3549 11491 -3545
rect 11427 -3605 11431 -3549
rect 11431 -3605 11487 -3549
rect 11487 -3605 11491 -3549
rect 11427 -3609 11491 -3605
rect 12595 -3549 12659 -3545
rect 12595 -3605 12599 -3549
rect 12599 -3605 12655 -3549
rect 12655 -3605 12659 -3549
rect 12595 -3609 12659 -3605
rect 13763 -3549 13827 -3545
rect 13763 -3605 13767 -3549
rect 13767 -3605 13823 -3549
rect 13823 -3605 13827 -3549
rect 13763 -3609 13827 -3605
rect 14931 -3549 14995 -3545
rect 14931 -3605 14935 -3549
rect 14935 -3605 14991 -3549
rect 14991 -3605 14995 -3549
rect 14931 -3609 14995 -3605
<< metal4 >>
rect 9865 1457 9931 1458
rect 9865 1393 9866 1457
rect 9930 1393 9931 1457
rect 9865 1392 9931 1393
rect 10419 1457 10485 1458
rect 10419 1393 10420 1457
rect 10484 1393 10485 1457
rect 10419 1392 10485 1393
rect 11113 1457 11179 1458
rect 11113 1393 11114 1457
rect 11178 1393 11179 1457
rect 11113 1392 11179 1393
rect 11667 1457 11733 1458
rect 11667 1393 11668 1457
rect 11732 1393 11733 1457
rect 11667 1392 11733 1393
rect 12361 1457 12427 1458
rect 12361 1393 12362 1457
rect 12426 1393 12427 1457
rect 12361 1392 12427 1393
rect 12915 1457 12981 1458
rect 12915 1393 12916 1457
rect 12980 1393 12981 1457
rect 12915 1392 12981 1393
rect 13609 1457 13675 1458
rect 13609 1393 13610 1457
rect 13674 1393 13675 1457
rect 13609 1392 13675 1393
rect 14163 1457 14229 1458
rect 14163 1393 14164 1457
rect 14228 1393 14229 1457
rect 14163 1392 14229 1393
rect 9580 337 9646 338
rect 9580 273 9581 337
rect 9645 273 9646 337
rect 9580 272 9646 273
rect 9090 -452 9156 -451
rect 9090 -516 9091 -452
rect 9155 -516 9156 -452
rect 9090 -517 9156 -516
rect 7922 -696 7988 -695
rect 7922 -760 7923 -696
rect 7987 -760 7988 -696
rect 7922 -761 7988 -760
rect 6754 -940 6820 -939
rect 6754 -1004 6755 -940
rect 6819 -1004 6820 -940
rect 6754 -1005 6820 -1004
rect 5586 -1184 5652 -1183
rect 5586 -1248 5587 -1184
rect 5651 -1248 5652 -1184
rect 5586 -1249 5652 -1248
rect 4418 -1428 4484 -1427
rect 4418 -1492 4419 -1428
rect 4483 -1492 4484 -1428
rect 4418 -1493 4484 -1492
rect 3250 -1672 3316 -1671
rect 3250 -1736 3251 -1672
rect 3315 -1736 3316 -1672
rect 3250 -1737 3316 -1736
rect 2082 -1916 2148 -1915
rect 2082 -1980 2083 -1916
rect 2147 -1980 2148 -1916
rect 2082 -1981 2148 -1980
rect 2085 -3544 2145 -1981
rect 3253 -3544 3313 -1737
rect 4421 -3544 4481 -1493
rect 5589 -3544 5649 -1249
rect 6757 -3544 6817 -1005
rect 7925 -3544 7985 -761
rect 9093 -3544 9153 -517
rect 9583 -1915 9643 272
rect 9868 -939 9928 1392
rect 10422 -695 10482 1392
rect 10828 337 10894 338
rect 10828 273 10829 337
rect 10893 273 10894 337
rect 10828 272 10894 273
rect 10419 -696 10485 -695
rect 10419 -760 10420 -696
rect 10484 -760 10485 -696
rect 10419 -761 10485 -760
rect 9865 -940 9931 -939
rect 9865 -1004 9866 -940
rect 9930 -1004 9931 -940
rect 9865 -1005 9931 -1004
rect 10258 -940 10324 -939
rect 10258 -1004 10259 -940
rect 10323 -1004 10324 -940
rect 10258 -1005 10324 -1004
rect 9580 -1916 9646 -1915
rect 9580 -1980 9581 -1916
rect 9645 -1980 9646 -1916
rect 9580 -1981 9646 -1980
rect 10261 -3544 10321 -1005
rect 10831 -1671 10891 272
rect 11116 -451 11176 1392
rect 11113 -452 11179 -451
rect 11113 -516 11114 -452
rect 11178 -516 11179 -452
rect 11113 -517 11179 -516
rect 11670 -939 11730 1392
rect 12076 337 12142 338
rect 12076 273 12077 337
rect 12141 273 12142 337
rect 12076 272 12142 273
rect 11667 -940 11733 -939
rect 11667 -1004 11668 -940
rect 11732 -1004 11733 -940
rect 11667 -1005 11733 -1004
rect 12079 -1427 12139 272
rect 12076 -1428 12142 -1427
rect 12076 -1492 12077 -1428
rect 12141 -1492 12142 -1428
rect 12076 -1493 12142 -1492
rect 12364 -1671 12424 1392
rect 10828 -1672 10894 -1671
rect 10828 -1736 10829 -1672
rect 10893 -1736 10894 -1672
rect 10828 -1737 10894 -1736
rect 11426 -1672 11492 -1671
rect 11426 -1736 11427 -1672
rect 11491 -1736 11492 -1672
rect 11426 -1737 11492 -1736
rect 12361 -1672 12427 -1671
rect 12361 -1736 12362 -1672
rect 12426 -1736 12427 -1672
rect 12361 -1737 12427 -1736
rect 11429 -3544 11489 -1737
rect 12918 -1915 12978 1392
rect 13324 337 13390 338
rect 13324 273 13325 337
rect 13389 273 13390 337
rect 13324 272 13390 273
rect 13327 -1183 13387 272
rect 13324 -1184 13390 -1183
rect 13324 -1248 13325 -1184
rect 13389 -1248 13390 -1184
rect 13324 -1249 13390 -1248
rect 13612 -1915 13672 1392
rect 14166 -1915 14226 1392
rect 12594 -1916 12660 -1915
rect 12594 -1980 12595 -1916
rect 12659 -1980 12660 -1916
rect 12594 -1981 12660 -1980
rect 12915 -1916 12981 -1915
rect 12915 -1980 12916 -1916
rect 12980 -1980 12981 -1916
rect 12915 -1981 12981 -1980
rect 13609 -1916 13675 -1915
rect 13609 -1980 13610 -1916
rect 13674 -1980 13675 -1916
rect 13609 -1981 13675 -1980
rect 13762 -1916 13828 -1915
rect 13762 -1980 13763 -1916
rect 13827 -1980 13828 -1916
rect 13762 -1981 13828 -1980
rect 14163 -1916 14229 -1915
rect 14163 -1980 14164 -1916
rect 14228 -1980 14229 -1916
rect 14163 -1981 14229 -1980
rect 14930 -1916 14996 -1915
rect 14930 -1980 14931 -1916
rect 14995 -1980 14996 -1916
rect 14930 -1981 14996 -1980
rect 12597 -3544 12657 -1981
rect 13765 -3544 13825 -1981
rect 14933 -3544 14993 -1981
rect 2082 -3545 2148 -3544
rect 2082 -3609 2083 -3545
rect 2147 -3609 2148 -3545
rect 2082 -3610 2148 -3609
rect 3250 -3545 3316 -3544
rect 3250 -3609 3251 -3545
rect 3315 -3609 3316 -3545
rect 3250 -3610 3316 -3609
rect 4418 -3545 4484 -3544
rect 4418 -3609 4419 -3545
rect 4483 -3609 4484 -3545
rect 4418 -3610 4484 -3609
rect 5586 -3545 5652 -3544
rect 5586 -3609 5587 -3545
rect 5651 -3609 5652 -3545
rect 5586 -3610 5652 -3609
rect 6754 -3545 6820 -3544
rect 6754 -3609 6755 -3545
rect 6819 -3609 6820 -3545
rect 6754 -3610 6820 -3609
rect 7922 -3545 7988 -3544
rect 7922 -3609 7923 -3545
rect 7987 -3609 7988 -3545
rect 7922 -3610 7988 -3609
rect 9090 -3545 9156 -3544
rect 9090 -3609 9091 -3545
rect 9155 -3609 9156 -3545
rect 9090 -3610 9156 -3609
rect 10258 -3545 10324 -3544
rect 10258 -3609 10259 -3545
rect 10323 -3609 10324 -3545
rect 10258 -3610 10324 -3609
rect 11426 -3545 11492 -3544
rect 11426 -3609 11427 -3545
rect 11491 -3609 11492 -3545
rect 11426 -3610 11492 -3609
rect 12594 -3545 12660 -3544
rect 12594 -3609 12595 -3545
rect 12659 -3609 12660 -3545
rect 12594 -3610 12660 -3609
rect 13762 -3545 13828 -3544
rect 13762 -3609 13763 -3545
rect 13827 -3609 13828 -3545
rect 13762 -3610 13828 -3609
rect 14930 -3545 14996 -3544
rect 14930 -3609 14931 -3545
rect 14995 -3609 14996 -3545
rect 14930 -3610 14996 -3609
use contact_30  contact_30_0
timestamp 1634918361
transform 1 0 9085 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1634918361
transform 1 0 9090 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_1
timestamp 1634918361
transform 1 0 9085 0 1 -517
box 0 0 1 1
use contact_30  contact_30_2
timestamp 1634918361
transform 1 0 11108 0 1 1392
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1634918361
transform 1 0 11113 0 1 1388
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1634918361
transform 1 0 11114 0 1 1393
box 0 0 1 1
use contact_30  contact_30_3
timestamp 1634918361
transform 1 0 11108 0 1 -517
box 0 0 1 1
use contact_30  contact_30_4
timestamp 1634918361
transform 1 0 7917 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1634918361
transform 1 0 7922 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_5
timestamp 1634918361
transform 1 0 7917 0 1 -761
box 0 0 1 1
use contact_30  contact_30_6
timestamp 1634918361
transform 1 0 10414 0 1 1392
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1634918361
transform 1 0 10419 0 1 1388
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1634918361
transform 1 0 10420 0 1 1393
box 0 0 1 1
use contact_30  contact_30_7
timestamp 1634918361
transform 1 0 10414 0 1 -761
box 0 0 1 1
use contact_30  contact_30_8
timestamp 1634918361
transform 1 0 10253 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1634918361
transform 1 0 10258 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_9
timestamp 1634918361
transform 1 0 10253 0 1 -1005
box 0 0 1 1
use contact_30  contact_30_10
timestamp 1634918361
transform 1 0 11662 0 1 1392
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1634918361
transform 1 0 11667 0 1 1388
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1634918361
transform 1 0 11668 0 1 1393
box 0 0 1 1
use contact_30  contact_30_11
timestamp 1634918361
transform 1 0 11662 0 1 -1005
box 0 0 1 1
use contact_30  contact_30_12
timestamp 1634918361
transform 1 0 6749 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1634918361
transform 1 0 6754 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_13
timestamp 1634918361
transform 1 0 6749 0 1 -1005
box 0 0 1 1
use contact_30  contact_30_14
timestamp 1634918361
transform 1 0 9860 0 1 1392
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1634918361
transform 1 0 9865 0 1 1388
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1634918361
transform 1 0 9866 0 1 1393
box 0 0 1 1
use contact_30  contact_30_15
timestamp 1634918361
transform 1 0 9860 0 1 -1005
box 0 0 1 1
use contact_30  contact_30_16
timestamp 1634918361
transform 1 0 5581 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1634918361
transform 1 0 5586 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_17
timestamp 1634918361
transform 1 0 5581 0 1 -1249
box 0 0 1 1
use contact_30  contact_30_18
timestamp 1634918361
transform 1 0 13319 0 1 272
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1634918361
transform 1 0 13324 0 1 268
box 0 0 1 1
use contact_30  contact_30_19
timestamp 1634918361
transform 1 0 13319 0 1 -1249
box 0 0 1 1
use contact_30  contact_30_20
timestamp 1634918361
transform 1 0 4413 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1634918361
transform 1 0 4418 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_21
timestamp 1634918361
transform 1 0 4413 0 1 -1493
box 0 0 1 1
use contact_30  contact_30_22
timestamp 1634918361
transform 1 0 12071 0 1 272
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1634918361
transform 1 0 12076 0 1 268
box 0 0 1 1
use contact_30  contact_30_23
timestamp 1634918361
transform 1 0 12071 0 1 -1493
box 0 0 1 1
use contact_30  contact_30_24
timestamp 1634918361
transform 1 0 11421 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1634918361
transform 1 0 11426 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_25
timestamp 1634918361
transform 1 0 11421 0 1 -1737
box 0 0 1 1
use contact_30  contact_30_26
timestamp 1634918361
transform 1 0 12356 0 1 1392
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1634918361
transform 1 0 12361 0 1 1388
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1634918361
transform 1 0 12362 0 1 1393
box 0 0 1 1
use contact_30  contact_30_27
timestamp 1634918361
transform 1 0 12356 0 1 -1737
box 0 0 1 1
use contact_30  contact_30_28
timestamp 1634918361
transform 1 0 3245 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1634918361
transform 1 0 3250 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_29
timestamp 1634918361
transform 1 0 3245 0 1 -1737
box 0 0 1 1
use contact_30  contact_30_30
timestamp 1634918361
transform 1 0 10823 0 1 272
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1634918361
transform 1 0 10828 0 1 268
box 0 0 1 1
use contact_30  contact_30_31
timestamp 1634918361
transform 1 0 10823 0 1 -1737
box 0 0 1 1
use contact_30  contact_30_32
timestamp 1634918361
transform 1 0 14925 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1634918361
transform 1 0 14930 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_33
timestamp 1634918361
transform 1 0 14925 0 1 -1981
box 0 0 1 1
use contact_30  contact_30_34
timestamp 1634918361
transform 1 0 14158 0 1 1392
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1634918361
transform 1 0 14163 0 1 1388
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1634918361
transform 1 0 14164 0 1 1393
box 0 0 1 1
use contact_30  contact_30_35
timestamp 1634918361
transform 1 0 14158 0 1 -1981
box 0 0 1 1
use contact_30  contact_30_36
timestamp 1634918361
transform 1 0 13757 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1634918361
transform 1 0 13762 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_37
timestamp 1634918361
transform 1 0 13757 0 1 -1981
box 0 0 1 1
use contact_30  contact_30_38
timestamp 1634918361
transform 1 0 13604 0 1 1392
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1634918361
transform 1 0 13609 0 1 1388
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1634918361
transform 1 0 13610 0 1 1393
box 0 0 1 1
use contact_30  contact_30_39
timestamp 1634918361
transform 1 0 13604 0 1 -1981
box 0 0 1 1
use contact_30  contact_30_40
timestamp 1634918361
transform 1 0 12589 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1634918361
transform 1 0 12594 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_41
timestamp 1634918361
transform 1 0 12589 0 1 -1981
box 0 0 1 1
use contact_30  contact_30_42
timestamp 1634918361
transform 1 0 12910 0 1 1392
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1634918361
transform 1 0 12915 0 1 1388
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1634918361
transform 1 0 12916 0 1 1393
box 0 0 1 1
use contact_30  contact_30_43
timestamp 1634918361
transform 1 0 12910 0 1 -1981
box 0 0 1 1
use contact_30  contact_30_44
timestamp 1634918361
transform 1 0 2077 0 1 -3610
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1634918361
transform 1 0 2082 0 1 -3614
box 0 0 1 1
use contact_30  contact_30_45
timestamp 1634918361
transform 1 0 2077 0 1 -1981
box 0 0 1 1
use contact_30  contact_30_46
timestamp 1634918361
transform 1 0 9575 0 1 272
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1634918361
transform 1 0 9580 0 1 268
box 0 0 1 1
use contact_30  contact_30_47
timestamp 1634918361
transform 1 0 9575 0 1 -1981
box 0 0 1 1
<< properties >>
string FIXED_BBOX 2040 -3614 15038 1462
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 1237220
string GDS_START 1229536
<< end >>
