magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1296 -1277 2042 2437
<< locali >>
rect 0 1103 746 1137
rect 212 485 246 551
rect 330 539 364 857
rect 330 505 459 539
rect 557 505 591 539
rect 112 237 146 303
rect 0 -17 746 17
use pdriver  pdriver_0
timestamp 1634918361
transform 1 0 378 0 1 0
box -36 -17 404 1177
use pnand2  pnand2_0
timestamp 1634918361
transform 1 0 0 0 1 0
box -36 -17 414 1177
<< labels >>
rlabel locali s 574 522 574 522 4 Z
port 1 nsew
rlabel locali s 129 270 129 270 4 A
port 2 nsew
rlabel locali s 229 518 229 518 4 B
port 3 nsew
rlabel locali s 373 0 373 0 4 gnd
port 4 nsew
rlabel locali s 373 1120 373 1120 4 vdd
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 746 1120
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 875350
string GDS_START 874280
<< end >>
