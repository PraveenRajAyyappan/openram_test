magic
tech sky130A
magscale 1 2
timestamp 1634918361
<< checkpaint >>
rect -1286 -1286 1436 1358
<< pwell >>
rect -26 -26 176 98
<< scnmos >>
rect 60 0 90 72
<< ndiff >>
rect 0 53 60 72
rect 0 19 8 53
rect 42 19 60 53
rect 0 0 60 19
rect 90 53 150 72
rect 90 19 108 53
rect 142 19 150 53
rect 90 0 150 19
<< ndiffc >>
rect 8 19 42 53
rect 108 19 142 53
<< poly >>
rect 60 72 90 98
rect 60 -26 90 0
<< locali >>
rect 8 53 42 69
rect 8 3 42 19
rect 108 53 142 69
rect 108 3 142 19
use contact_11  contact_11_0
timestamp 1634918361
transform 1 0 100 0 1 3
box 0 0 1 1
use contact_11  contact_11_1
timestamp 1634918361
transform 1 0 0 0 1 3
box 0 0 1 1
<< labels >>
rlabel poly s 75 36 75 36 4 G
port 1 nsew
rlabel locali s 25 36 25 36 4 S
port 2 nsew
rlabel locali s 125 36 125 36 4 D
port 3 nsew
<< properties >>
string FIXED_BBOX -25 -26 175 98
string GDS_FILE sky130_sram_0kbytes_1rw1r_8x16_2.gds
string GDS_END 884682
string GDS_START 883954
<< end >>
